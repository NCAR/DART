netcdf filter_input {
dimensions:
	member = 20 ;
	metadatalength = 32 ;
	location = 9 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;

	double state(time, member, location) ;
		state:long_name = "the ensemble of model states" ;

	double state_priorinf_mean(time, location) ;
		state_priorinf_mean:long_name = "prior inflation value" ;

	double state_priorinf_sd(time, location) ;
		state_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double state_postinf_mean(time, location) ;
		state_postinf_mean:long_name = "posterior inflation value" ;

	double state_postinf_sd(time, location) ;
		state_postinf_sd:long_name = "posterior inflation standard deviation" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "days" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
                :model = "9var" ;
                :model_g = 8. ;
                :model_deltat = 0.0833333333333333 ;
                :model_a = 1., 1., 3. ;
                :model_b = -1.5, -1.5, 0.5 ;
                :model_f = 0.1, 0., 0. ;
                :model_h = -1., 0., 0. ;
                :model_nu = 0.0208333333333333 ;
                :model_kappa = 0.0208333333333333 ;
                :model_c = 0.8660254 ;
		:history = "identical (within 64bit precision) to filter_ics r1330 (circa June 2005)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20" ;

 location = 0, 0.111111111111111, 0.222222222222222, 0.333333333333333,
    0.444444444444444, 0.555555555555556, 0.666666666666667,
    0.777777777777778, 0.888888888888889 ;

 state =
 -1.106862221544870E-002, 3.771290104870961E-003, -4.267924910635314E-004,
    0.114948589376236     , -4.675421446496910E-003, -3.144985685982593E-002,
    0.114771987522227     , 3.315034128905045E-004, -3.103789754682037E-002,
 -1.097629908544451E-002, 1.628870120884410E-003, -1.724367100664169E-003,
    0.153884898469423     , -4.609178488475665E-002, -1.074826135017564E-002,
    0.153376419620458     , -4.353771179526299E-002, -7.330011764484777E-003,
 -1.115601895285006E-002, -2.121639701918137E-003, -3.663403642228576E-004,
    0.184167211396182     , -1.565068707325053E-002, 1.685168248189148E-002,
    0.184738134390312     , -2.004376155667765E-002, 1.810159492670806E-002,
 -1.151689848629175E-002, -8.172881282684098E-003, 2.140196049682653E-005,
 -6.498925306326872E-002, -1.469979932167828E-002, 9.610790680442356E-002,
 -6.444693139132428E-002, -3.358379026676453E-003, 9.517561713228902E-002,
 -1.115703091688085E-002, -2.414458777888068E-003, -2.916829013787560E-004,
    0.171419940206066     , -1.400123030376602E-002, 1.932706155775381E-002,
    0.171983781722834     , -1.867949404070250E-002, 2.033285515268970E-002,
 -1.101477765809463E-002, -4.739645804187219E-003, 6.470948260225287E-004,
    8.345520919944314E-002, 9.666897541339299E-003, 4.133314427015217E-002,
    8.276304634271292E-002, 5.069681705867740E-003, 4.078700726980420E-002,
 -1.112284391099167E-002, 1.984844657211081E-003, 2.473035703491002E-005,
    0.179073062377889     , 5.415261119287277E-003, -1.543651481109227E-002,
    0.179383687146613     , 9.360359734681231E-003, -1.578670996051275E-002,
 -1.097910442221214E-002, 1.517238090950208E-003, -1.789099020026624E-003,
    0.155514522823682     , -4.819161259442939E-002, -9.738341108145563E-003,
    0.155050458810241     , -4.582384708692750E-002, -6.133882290120902E-003,
 -1.113275521794145E-002, 2.294332251740906E-003, 8.402898535670641E-005,
    0.170164019681455     , 7.727169238560596E-003, -1.813345989946173E-002,
    0.170541591185717     , 1.210655078009050E-002, -1.863258552349303E-002,
 -1.109935551170690E-002, 1.447728648448185E-003, -2.547946512265806E-004,
    0.189540824861343     , -3.819823837293403E-003, -1.073482194562231E-002,
    0.189689904960803     , -8.673372379088949E-004, -1.030665950805344E-002,
 -1.071841648321390E-002, -5.900078717788844E-003, 1.544266608899803E-003,
    4.323479035823961E-002, 3.406523598464715E-002, 5.373094717557179E-002,
    4.018369001215370E-002, 3.131559684765405E-002, 5.293890489406514E-002,
 -1.447465875170160E-002, -8.202008235743043E-003, -9.047052148967812E-003,
    0.143966427509255     , -0.264683263240974     , 8.068344281367744E-002,
    0.175464380438600     , -0.279804742835901     , 9.776963982259521E-002,
 -1.098608930470730E-002, 1.563594455526852E-003, -1.666148933613321E-003,
    0.156184109229457     , -4.453803377826222E-002, -1.026421981433804E-002,
    0.155733316460666     , -4.205966467049859E-002, -6.909847867764780E-003,
 -1.116422244942031E-002, -2.319082215120003E-003, -3.896542413340770E-004,
    0.177528006128431     , -1.669191241809743E-002, 1.856364203489457E-002,
    0.178156209767679     , -2.134448410032458E-002, 1.984106768608409E-002,
 -1.107830651013313E-002, 1.055708749500965E-003, -7.023719749990172E-004,
    0.189479321879420     , -1.768969803408101E-002, -7.129031617637074E-003,
    0.189516926295396     , -1.565805212094398E-002, -5.472307194241021E-003,
 -1.079096822101823E-002, -4.683208804437237E-003, 1.556441399616348E-003,
    8.025690201240224E-002, 3.607802754049073E-002, 3.967889907664456E-002,
    7.806196154000131E-002, 3.174850029013718E-002, 3.821318691268807E-002,
 -1.110832336062493E-002, -3.547645027200915E-003, 2.044743315014535E-004,
    0.125370868974225     , -1.443023385685434E-003, 2.940167067707648E-002,
    0.125500172663210     , -6.569349739277322E-003, 2.932435333843108E-002,
 -1.489761967487414E-002, -8.381405068944591E-003, -6.090343246197891E-003,
   -2.185857229057468E-002, -0.181405371959135     , 0.104393803185557     ,
    4.987290816873804E-003, -0.175311586925613     , 0.100689174193223     ,
 -1.111955578092320E-002, 3.231517899165453E-003, -1.174403580331110E-004,
    0.135993377636909     , 3.466525655903596E-003, -2.646283904792186E-002,
    0.136227689279231     , 8.502730383204071E-003, -2.653006786332830E-002,
 -1.112043735652409E-002, -1.642273506646009E-003, -4.095338601362411E-005,
    0.191822867067069     , -5.209167449539595E-003, 1.258790297239439E-002,
    0.192121871082892     , -8.669700488602243E-003, 1.296840222515883E-002 ;

 state_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 state_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 state_postinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 state_postinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 time = 249.75 ;

 advance_to_time = 249.75 ;
}
