netcdf filter_input_source_noise {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 10 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double concentration(time, member, location) ;
		concentration:long_name = "tracer concentration" ;
		concentration:units = "mass" ;

	double mean_source(time, member, location) ;
		mean_source:long_name = "mean source" ;
		mean_source:units = "mass/timestep" ;

	double source(time, member, location) ;
		source:long_name = "source" ;
		source:units = "mass/timestep" ;

	double source_phase(time, member, location) ;
		source_phase:long_name = "source phase" ;
		source_phase:units = "radians" ;

	double wind(time, member, location) ;
		wind:long_name = "wind" ;
		wind:units = "gridpoints/timestep" ;

	double concentration_priorinf_mean(time, location) ;
		concentration_priorinf_mean:long_name = "prior inflation value for concentration" ;

	double mean_source_priorinf_mean(time, location) ;
		mean_source_priorinf_mean:long_name = "prior inflation value for mean source" ;

	double source_phase_priorinf_mean(time, location) ;
		source_phase_priorinf_mean:long_name = "prior inflation value for source phase" ;

	double source_priorinf_mean(time, location) ;
		source_priorinf_mean:long_name = "prior inflation value for source" ;

	double wind_priorinf_mean(time, location) ;
		wind_priorinf_mean:long_name = "prior inflation value for wind" ;

	double concentration_priorinf_sd(time, location) ;
		concentration_priorinf_sd:long_name = "prior inflation standard deviation for concentration" ;

	double mean_source_priorinf_sd(time, location) ;
		mean_source_priorinf_sd:long_name = "prior inflation standard deviation for mean source" ;

	double source_phase_priorinf_sd(time, location) ;
		source_phase_priorinf_sd:long_name = "prior inflation standard deviation for source phase" ;

	double source_priorinf_sd(time, location) ;
		source_priorinf_sd:long_name = "prior inflation standard deviation for source" ;

	double wind_priorinf_sd(time, location) ;
		wind_priorinf_sd:long_name = "prior inflation standard deviation for wind" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;
		location:axis = "X" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "days" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
                :description = "Initial conditions for varying source model experiments." ; 
		:model = "simple_advection" ;
		:destruction_rate = 5.555556e-05 ;
		:history = "same values as in filter_ics r3004 (circa July 2007)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 concentration =
  4894.89912670214, 4105.75196046983, 3300.69425212921, 2859.2620617744, 
    2539.94023370335, 2205.44300854388, 2054.83918208125, 1903.71154654458, 
    1753.33322606873, 1677.23096004728,
  4790.16331006911, 4122.07548155903, 3356.48669022321, 2841.52592353415, 
    2534.67990171862, 2221.88714285059, 2090.01851075256, 1892.9305518882, 
    1742.63612902049, 1699.3026495544,
  4880.78033245294, 4117.5511649177, 3313.53703565025, 2903.9950388971, 
    2510.20725030002, 2215.95689428705, 2058.48181442404, 1873.73221059902, 
    1723.10156995026, 1685.12867561787,
  4848.65398467122, 4137.48584245974, 3291.68069595039, 2849.9503014071, 
    2541.50696380899, 2286.78532017773, 2078.31316876191, 1874.02192423749, 
    1766.08267232634, 1674.70342488489,
  4937.0929593071, 4026.34481600101, 3327.7571275614, 2914.68740102219, 
    2632.55772487232, 2253.15521200829, 2058.97684997662, 1906.55469689961, 
    1741.31332898544, 1684.7526694428,
  4790.82174879002, 4006.27728404875, 3325.62332918537, 2930.42934958294, 
    2528.93815261724, 2223.94445225081, 2027.61432746, 1854.45138323444, 
    1742.93980770942, 1660.22383962852,
  4847.97907517179, 4096.1802838888, 3365.81551867447, 2860.4504863709, 
    2538.2512425897, 2235.73201597637, 2043.92469427129, 1914.90783158837, 
    1734.42565449291, 1669.52439435519,
  4914.04241591443, 4076.80309900796, 3301.00676933442, 2847.75024048709, 
    2486.84037046482, 2218.89171525289, 2064.22609372495, 1891.06190675184, 
    1771.75632681588, 1679.28947495859,
  4881.62237436124, 4046.85673163887, 3370.44473310472, 2868.19633695997, 
    2542.14297840282, 2204.75689059446, 2096.75964541014, 1908.97639278675, 
    1748.15389161777, 1666.13990112217,
  4762.58297087179, 4049.38410784739, 3382.48169841102, 2858.81153566859, 
    2500.80072574183, 2216.07192309216, 2031.95679693811, 1899.01836943805, 
    1763.39090540807, 1654.99953593773,
  4870.10979755572, 4060.08004860176, 3288.42095219066, 2864.95843791304, 
    2509.46934125534, 2239.47647952268, 2082.72036095693, 1911.06004631412, 
    1748.22786671053, 1649.82345814584,
  4857.13543681385, 4116.5327689139, 3333.27666106003, 2908.53154631149, 
    2528.12578319159, 2207.43608189493, 2024.65311280384, 1916.37387209997, 
    1727.83818240331, 1665.93182864471,
  4837.26234542043, 4088.74282516886, 3330.47337717606, 2886.17299193205, 
    2539.6105773162, 2234.09827101964, 2049.63623696516, 1891.96446908575, 
    1737.23160707505, 1689.85233045729,
  4888.62678243545, 4030.73870664674, 3338.81583537355, 2880.77658203231, 
    2493.10299066874, 2278.32391110113, 2055.47171724203, 1870.1588276368, 
    1760.51842798513, 1651.94992035752,
  4851.84811189662, 4128.45875046487, 3314.44264662302, 2948.20147280166, 
    2481.98207304599, 2249.87570743147, 2048.87979530252, 1872.88851346332, 
    1790.70602169075, 1673.06190920683,
  4878.25425690904, 4099.14890560483, 3303.01809989407, 2920.23892741273, 
    2514.534654533, 2222.47598907938, 2038.86022582934, 1891.17784986293, 
    1746.50212752721, 1680.52838298128,
  4890.04290777119, 4078.27426695272, 3377.76158625823, 2875.76601973321, 
    2548.32068016111, 2223.45994590661, 2041.20619064588, 1930.1812180781, 
    1769.39393988508, 1680.225276927,
  4784.92528667434, 4093.79062483647, 3280.60629651322, 2834.74218300042, 
    2524.66790706486, 2228.33598639446, 2045.74691644795, 1893.31506518768, 
    1739.55935925178, 1693.71272828427,
  4805.47251863082, 4107.68272480209, 3297.53762046689, 2872.67479263842, 
    2554.39660255678, 2229.35114248145, 2066.0945609762, 1878.40426522738, 
    1741.50209547843, 1672.36456265195,
  4857.56878063194, 4082.81870133308, 3399.89871220814, 2850.28266865423, 
    2572.57622489846, 2250.17592997059, 2029.23096607576, 1876.27664855374, 
    1761.99618821085, 1683.31669846937,
  4897.28261228406, 4049.5200161417, 3333.24340755026, 2868.76368054753, 
    2544.09412810106, 2242.05294119562, 2051.70230807087, 1883.61717148667, 
    1706.89822653913, 1658.95811711011,
  4886.04441292312, 4054.56002893158, 3314.63349048205, 2904.91436425581, 
    2497.66955442718, 2258.19536598303, 2061.57034789758, 1885.6897383932, 
    1743.34780226748, 1675.78018190345,
  4766.70342911952, 4126.81116891038, 3321.12728430556, 2899.08422025579, 
    2553.02927045044, 2212.66156303798, 2044.99309725918, 1905.16972544504, 
    1745.8982454938, 1665.54247405791,
  4810.76134560102, 4057.24825065536, 3388.20214667225, 2792.20640318031, 
    2534.65416269188, 2249.43615453335, 2026.82403030901, 1876.7455071391, 
    1759.58124628428, 1691.35495285619,
  4800.42074511709, 4083.36744442034, 3308.64120538478, 2879.35079154502, 
    2532.40593509346, 2264.31401438522, 2047.43236889578, 1884.45408951449, 
    1749.2138006992, 1681.35903947328,
  4821.36674841851, 4116.44364885516, 3316.65559651036, 2866.08708914746, 
    2542.55825472408, 2229.00052588989, 2048.28589832738, 1891.32231537889, 
    1774.30534229716, 1717.81240371683,
  4877.39528435894, 4043.80932351187, 3339.17470264656, 2862.17389234546, 
    2502.98882665194, 2234.72100156208, 2036.86625174707, 1897.86743187548, 
    1779.22266696005, 1700.41266308539,
  4825.48704294234, 4066.02924798193, 3286.64300346579, 2939.26783478542, 
    2541.99224376877, 2220.75760221135, 2021.02582710213, 1906.67803714594, 
    1749.70173828488, 1692.6833335697,
  4843.70313539504, 4065.13832690927, 3301.05445011417, 2882.03903897785, 
    2568.47078408025, 2211.12859016757, 2048.03849074765, 1864.39023874517, 
    1749.96974079079, 1666.57936469885,
  4872.48475495851, 4064.33945014901, 3342.2144591961, 2866.62298543211, 
    2553.20311298233, 2247.71883013158, 2046.09146519222, 1914.42032750192, 
    1772.69129574734, 1669.86264975504,
  4768.70766373274, 4052.50739436061, 3300.96718967926, 2901.79371862174, 
    2519.70681530917, 2227.86683132498, 2047.12325310543, 1905.64469415517, 
    1750.99082419178, 1683.72528475088,
  4794.90316947322, 4128.64405340403, 3313.65657469427, 2856.56948078172, 
    2572.96269258333, 2261.29545640129, 2046.4150204607, 1884.68240417412, 
    1782.21888699291, 1698.70022377959,
  4861.14020632389, 3963.96419873824, 3311.23023438765, 2830.87529624295, 
    2538.97267444093, 2203.1874367338, 2083.36879799288, 1891.69794173375, 
    1751.47450942309, 1692.21462619422,
  4798.54811625812, 4070.68304439599, 3288.53853386342, 2879.33676180386, 
    2505.4432295262, 2256.85431681328, 2057.093777098, 1881.06515769021, 
    1745.64887835977, 1683.74432385239,
  4842.91963620633, 4079.60020962004, 3335.53025316483, 2849.52259786707, 
    2524.68620965972, 2279.5720437524, 2049.15529077205, 1891.93212191096, 
    1751.02844517101, 1674.37440597125,
  4750.86022824831, 4087.0454315121, 3330.70205824596, 2832.0941765725, 
    2493.52534630975, 2226.84574629272, 2039.76766863019, 1893.25114275368, 
    1747.72981479267, 1679.04440397231,
  4810.13991926841, 4099.43563485646, 3355.89314980616, 2917.58359984831, 
    2522.58005394742, 2254.50231826997, 2035.00896127076, 1889.52336519947, 
    1760.94735130471, 1692.32733060092,
  4796.62587919365, 4084.34858686292, 3299.71397372026, 2852.5641914817, 
    2542.27941803384, 2263.56518698657, 2046.12646045433, 1899.86303878244, 
    1762.02634337594, 1695.69056503413,
  4885.79422130652, 4070.80571757784, 3367.93829038464, 2856.00866219034, 
    2517.16345003706, 2263.54200436205, 2021.16388006763, 1840.47882069779, 
    1756.24485845195, 1682.96019862892,
  4807.92975218382, 4085.34920598337, 3385.77326114449, 2896.10210634008, 
    2533.7880933302, 2209.59864237498, 2070.52402569892, 1881.43949883564, 
    1748.42927876495, 1678.65299904054,
  4838.29230237748, 4117.92467283603, 3391.31037463279, 2841.04151227149, 
    2549.76387414836, 2237.0520233191, 2056.60909602614, 1899.24379047321, 
    1728.27102696581, 1677.22483840766,
  4768.73139341517, 4101.29992068724, 3299.78562977923, 2874.19759570816, 
    2520.13958328409, 2261.31541198439, 2074.88314951981, 1899.70570633978, 
    1753.98308202598, 1687.08985607122,
  4823.29980979498, 4079.30977364043, 3312.59474684216, 2870.04306162814, 
    2587.24918243282, 2253.50529667011, 2043.63627207111, 1872.20938593059, 
    1748.38132950368, 1665.82644742571,
  4839.38038663675, 4063.09100055982, 3332.9205627305, 2869.23753905632, 
    2572.99262259474, 2210.53096563062, 2060.06702967432, 1869.43287415312, 
    1769.81107088735, 1679.51161267801,
  4857.65987317818, 4069.38666214629, 3336.99807213275, 2879.17041079465, 
    2515.77847940871, 2249.89508815996, 2055.24131389157, 1887.36540060167, 
    1749.31728640906, 1689.06224655817,
  4857.5906284953, 4077.20611700515, 3361.76198950585, 2856.29443823018, 
    2533.22622074157, 2208.92879086953, 2061.42766745061, 1896.85120062051, 
    1807.52854737915, 1685.54641736585,
  4905.98774853182, 4053.30208950418, 3260.83884290556, 2903.25074330157, 
    2490.5659921835, 2183.56642001064, 2033.86743172255, 1890.53936663663, 
    1718.12330635835, 1670.47979445963,
  4841.75855188679, 4074.72561909215, 3317.41727535708, 2854.84304894942, 
    2563.49983279056, 2246.06080574137, 2041.49873712799, 1872.94057411632, 
    1737.57102870412, 1661.54572081924,
  4827.23259838231, 4051.13782056697, 3301.99161376605, 2892.80786697589, 
    2509.11380713777, 2261.58045372737, 2081.88189112021, 1893.58059485513, 
    1758.51450109442, 1687.80871998161,
  4798.50773131575, 4133.43560668014, 3289.70358831435, 2884.48086762671, 
    2518.51810073314, 2208.21815490436, 2031.61119583154, 1902.37441088168, 
    1759.58506993277, 1693.29076211151,
  4856.77680774253, 4050.07423283141, 3292.11365173481, 2901.95153781962, 
    2567.47751117913, 2231.3043332988, 2035.69744172239, 1874.72371893234, 
    1762.23193891912, 1712.34980726265,
  4848.86237228298, 4048.31650003213, 3317.51283305729, 2864.97122926436, 
    2462.5448049424, 2259.66446967668, 2053.85630358089, 1888.13252087839, 
    1745.23206884758, 1676.81517439388,
  4862.41609298508, 4071.99182675966, 3324.2950437095, 2862.9780106374, 
    2487.28240663281, 2296.6911788747, 2046.16873508969, 1938.68450873113, 
    1744.94974108117, 1702.54639180138,
  4876.01221520061, 4055.5647448987, 3285.26478878713, 2878.68285679989, 
    2522.39196225615, 2231.09301423885, 1994.08999252312, 1907.99559472248, 
    1774.04518883897, 1683.0482464109,
  4792.17973275548, 4097.94244737828, 3361.54108010218, 2864.51803528892, 
    2522.2935415644, 2241.14052241558, 2079.0076339587, 1876.36008072074, 
    1743.27193078483, 1692.54696751931,
  4904.25744936242, 4077.16461977851, 3349.59798111034, 2888.36434806296, 
    2510.00329874125, 2217.31475022811, 2085.21264587599, 1901.58931033077, 
    1754.9566695765, 1679.23952679011,
  4840.20585886782, 4054.97924476707, 3340.14623114307, 2857.39925152742, 
    2524.32124161694, 2221.06715965344, 2017.00557810896, 1913.97899805584, 
    1733.92875044847, 1672.85381122751,
  4831.74909388443, 4108.57162304925, 3285.33935852964, 2916.69248002291, 
    2517.55211867603, 2260.63915563959, 2064.0864013317, 1871.18651539646, 
    1746.95999511155, 1684.44746622932,
  4809.09623617218, 4140.16314163765, 3317.29078306703, 2834.76509051723, 
    2511.40020016064, 2234.26185435351, 2054.25204015457, 1889.24938886097, 
    1758.09199699033, 1682.08984946201,
  4781.55334917222, 4082.81201216679, 3304.14592249908, 2863.53269012893, 
    2544.67511945714, 2231.38340252312, 2058.47415369053, 1882.35382969834, 
    1747.8821265338, 1674.20193273918,
  4834.01154169747, 4048.23034185939, 3403.57836602231, 2844.36534433393, 
    2562.38925847696, 2223.64675758416, 2054.56648339253, 1877.31317051713, 
    1748.02987221783, 1676.47541749847,
  4841.01974271912, 4058.57793110009, 3373.42174174812, 2918.83479770857, 
    2511.19148319057, 2242.5540788056, 2035.63084793734, 1869.82351746595, 
    1766.55619467829, 1674.13331778648,
  4928.96300408838, 4051.39060286015, 3341.55989859557, 2905.12387223258, 
    2497.65358722319, 2245.55935966636, 2058.91130481889, 1914.53961913824, 
    1744.1251737207, 1657.8874893352,
  4845.93928119666, 4053.98204310441, 3329.5353467599, 2811.52820676734, 
    2557.30158420434, 2263.5915110411, 2057.70305392287, 1897.7171229324, 
    1750.08528934515, 1663.96572166461,
  4789.69598810755, 4116.7258309323, 3337.35047500115, 2864.83120364006, 
    2527.58491294468, 2208.87217988188, 2032.96890891952, 1853.76667575728, 
    1731.59261980527, 1684.24239889101,
  4801.72382140507, 4030.79349187825, 3305.9946565004, 2887.85515433118, 
    2563.68693540893, 2193.8866797347, 2046.16222941391, 1925.79738309505, 
    1753.2269054008, 1684.30580328263,
  4934.3586411042, 4069.77532160807, 3304.89315827795, 2862.6140435541, 
    2549.77698301134, 2243.21744471985, 2068.36938000894, 1869.13784081027, 
    1749.60350607073, 1668.74343675644,
  4825.86693860514, 4092.75002777421, 3332.34201597937, 2902.8991228243, 
    2537.99360751218, 2220.5238904846, 2069.56801926602, 1875.88390153588, 
    1742.35546941336, 1681.51725967009,
  4806.52827128191, 4076.70092005298, 3290.480416807, 2927.29919195151, 
    2521.7459395147, 2240.21181385823, 2047.65989812636, 1876.4589969647, 
    1760.78154940062, 1695.09927252104,
  4710.14802963826, 4126.078398214, 3325.85970012827, 2963.78889166522, 
    2533.95228806005, 2249.90839096506, 2111.9363519683, 1904.94338607073, 
    1757.36812245237, 1695.63326347093,
  4768.23828597436, 4102.57422667745, 3355.15664805721, 2864.11810079416, 
    2534.48055204207, 2224.71586369144, 2056.00650801869, 1907.30242662277, 
    1750.31275712004, 1676.22379522444,
  4816.44329423605, 4041.39564491723, 3336.13387186639, 2824.32821799534, 
    2598.28756657445, 2250.99042162813, 2037.37096012798, 1866.6101759189, 
    1739.63710542033, 1678.30898426862,
  4882.93678586238, 4107.2771317462, 3296.88485480303, 2883.58298411646, 
    2561.94923388669, 2256.03554964951, 2059.39453025837, 1909.78255837806, 
    1750.79876789948, 1676.82534020295,
  4772.4527063711, 4127.47604864852, 3240.65274897576, 2897.75789052099, 
    2499.71526860494, 2267.22232737705, 2051.65051633163, 1898.92774275018, 
    1743.01511080737, 1690.46137982271,
  4898.38050255964, 4060.98186475414, 3318.96684053055, 2842.45657674031, 
    2558.16199052052, 2213.52431275024, 2028.84122087278, 1880.23010395246, 
    1761.18990387355, 1686.10329799372,
  4801.11670447972, 4071.28858658671, 3326.84643227664, 2850.67508615821, 
    2558.89848335376, 2258.78800244523, 2037.80901117458, 1939.81364621208, 
    1783.43840441455, 1670.03829062678,
  4920.49250212555, 4085.19574151074, 3310.79129919349, 2849.52852973404, 
    2551.70912175383, 2239.93604727114, 2045.4773256901, 1882.11431007984, 
    1748.86361886835, 1661.04050239777,
  4831.41753828055, 4100.0081376777, 3326.72503950126, 2878.59731095118, 
    2533.80461804525, 2232.93043719701, 2063.5378000473, 1919.1631457192, 
    1774.66232867102, 1682.27811183685,
  4829.54899269637, 4065.64638393322, 3344.43647527355, 2946.23454974271, 
    2523.79728795556, 2273.11025760936, 2036.51858902943, 1914.08052369881, 
    1766.73761529178, 1691.0405041948,
  4849.16421069555, 4047.47100427488, 3312.3120381535, 2876.32290598557, 
    2534.0176456632, 2202.42397239549, 2060.59312314399, 1891.60031477213, 
    1753.4270559813, 1701.11422830225 ;

 mean_source =
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.00000000000249, 0.100000000000248, 0.100000000000248, 0.100000000000248, 
    0.100000000000248, 0.100000000000248, 0.100000000000248, 
    0.100000000000248, 0.100000000000248, 0.100000000000248,
  1.00000000000242, 0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241,
  1.00000000000257, 0.100000000000256, 0.100000000000256, 0.100000000000256, 
    0.100000000000256, 0.100000000000256, 0.100000000000256, 
    0.100000000000256, 0.100000000000256, 0.100000000000256,
  1.00000000000262, 0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261,
  1.0000000000025, 0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249,
  1.00000000000244, 0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243,
  1.0000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025,
  1.00000000000264, 0.100000000000263, 0.100000000000263, 0.100000000000263, 
    0.100000000000263, 0.100000000000263, 0.100000000000263, 
    0.100000000000263, 0.100000000000263, 0.100000000000263,
  1.00000000000252, 0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251,
  1.00000000000249, 0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249,
  1.00000000000254, 0.100000000000253, 0.100000000000253, 0.100000000000253, 
    0.100000000000253, 0.100000000000253, 0.100000000000253, 
    0.100000000000253, 0.100000000000253, 0.100000000000253,
  1.00000000000246, 0.100000000000246, 0.100000000000246, 0.100000000000246, 
    0.100000000000246, 0.100000000000246, 0.100000000000246, 
    0.100000000000246, 0.100000000000246, 0.100000000000246,
  1.00000000000243, 0.100000000000242, 0.100000000000242, 0.100000000000242, 
    0.100000000000242, 0.100000000000242, 0.100000000000242, 
    0.100000000000242, 0.100000000000242, 0.100000000000242,
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.00000000000254, 0.100000000000253, 0.100000000000253, 0.100000000000253, 
    0.100000000000253, 0.100000000000253, 0.100000000000253, 
    0.100000000000253, 0.100000000000253, 0.100000000000253,
  1.00000000000251, 0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251,
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.0000000000024, 0.100000000000239, 0.100000000000239, 0.100000000000239, 
    0.100000000000239, 0.100000000000239, 0.100000000000239, 
    0.100000000000239, 0.100000000000239, 0.100000000000239,
  1.00000000000251, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025,
  1.00000000000246, 0.100000000000245, 0.100000000000245, 0.100000000000245, 
    0.100000000000245, 0.100000000000245, 0.100000000000245, 
    0.100000000000245, 0.100000000000245, 0.100000000000245,
  1.00000000000248, 0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247,
  1.00000000000252, 0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251,
  1.00000000000248, 0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247,
  1.00000000000236, 0.100000000000236, 0.100000000000236, 0.100000000000236, 
    0.100000000000236, 0.100000000000236, 0.100000000000236, 
    0.100000000000236, 0.100000000000236, 0.100000000000236,
  1.00000000000263, 0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262,
  1.00000000000244, 0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243,
  1.00000000000241, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024,
  1.0000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025,
  1.00000000000263, 0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262,
  1.00000000000255, 0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255,
  1.00000000000243, 0.100000000000242, 0.100000000000242, 0.100000000000242, 
    0.100000000000242, 0.100000000000242, 0.100000000000242, 
    0.100000000000242, 0.100000000000242, 0.100000000000242,
  1.00000000000258, 0.100000000000257, 0.100000000000257, 0.100000000000257, 
    0.100000000000257, 0.100000000000257, 0.100000000000257, 
    0.100000000000257, 0.100000000000257, 0.100000000000257,
  1.00000000000261, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026,
  1.00000000000255, 0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255,
  1.0000000000024, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024,
  1.00000000000256, 0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255,
  1.0000000000024, 0.100000000000239, 0.100000000000239, 0.100000000000239, 
    0.100000000000239, 0.100000000000239, 0.100000000000239, 
    0.100000000000239, 0.100000000000239, 0.100000000000239,
  1.00000000000248, 0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247,
  1.00000000000258, 0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258,
  1.00000000000262, 0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262, 
    0.100000000000262, 0.100000000000262, 0.100000000000262,
  1.00000000000251, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025,
  1.00000000000259, 0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258,
  1.00000000000242, 0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241,
  1.00000000000261, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026,
  1.00000000000248, 0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247,
  1.00000000000253, 0.100000000000252, 0.100000000000252, 0.100000000000252, 
    0.100000000000252, 0.100000000000252, 0.100000000000252, 
    0.100000000000252, 0.100000000000252, 0.100000000000252,
  1.00000000000255, 0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254,
  1.0000000000025, 0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249,
  1.00000000000241, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024, 0.10000000000024, 0.10000000000024, 
    0.10000000000024, 0.10000000000024,
  1.00000000000244, 0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243,
  1.00000000000262, 0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261,
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.00000000000252, 0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251, 
    0.100000000000251, 0.100000000000251, 0.100000000000251,
  1.00000000000236, 0.100000000000235, 0.100000000000235, 0.100000000000235, 
    0.100000000000235, 0.100000000000235, 0.100000000000235, 
    0.100000000000235, 0.100000000000235, 0.100000000000235,
  1.00000000000238, 0.100000000000237, 0.100000000000237, 0.100000000000237, 
    0.100000000000237, 0.100000000000237, 0.100000000000237, 
    0.100000000000237, 0.100000000000237, 0.100000000000237,
  1.00000000000253, 0.100000000000252, 0.100000000000252, 0.100000000000252, 
    0.100000000000252, 0.100000000000252, 0.100000000000252, 
    0.100000000000252, 0.100000000000252, 0.100000000000252,
  1.00000000000246, 0.100000000000245, 0.100000000000245, 0.100000000000245, 
    0.100000000000245, 0.100000000000245, 0.100000000000245, 
    0.100000000000245, 0.100000000000245, 0.100000000000245,
  1.00000000000261, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026, 0.10000000000026, 0.10000000000026, 
    0.10000000000026, 0.10000000000026,
  1.00000000000237, 0.100000000000237, 0.100000000000237, 0.100000000000237, 
    0.100000000000237, 0.100000000000237, 0.100000000000237, 
    0.100000000000237, 0.100000000000237, 0.100000000000237,
  1.00000000000259, 0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258,
  1.00000000000251, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025, 0.10000000000025, 0.10000000000025, 
    0.10000000000025, 0.10000000000025,
  1.00000000000254, 0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254,
  1.0000000000025, 0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249,
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.00000000000236, 0.100000000000235, 0.100000000000235, 0.100000000000235, 
    0.100000000000235, 0.100000000000235, 0.100000000000235, 
    0.100000000000235, 0.100000000000235, 0.100000000000235,
  1.00000000000244, 0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243, 
    0.100000000000243, 0.100000000000243, 0.100000000000243,
  1.00000000000255, 0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254,
  1.00000000000243, 0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241, 
    0.100000000000241, 0.100000000000241, 0.100000000000241,
  1.00000000000269, 0.100000000000268, 0.100000000000268, 0.100000000000268, 
    0.100000000000268, 0.100000000000268, 0.100000000000268, 
    0.100000000000268, 0.100000000000268, 0.100000000000268,
  1.00000000000258, 0.100000000000257, 0.100000000000257, 0.100000000000257, 
    0.100000000000257, 0.100000000000257, 0.100000000000257, 
    0.100000000000257, 0.100000000000257, 0.100000000000257,
  1.00000000000248, 0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247, 
    0.100000000000247, 0.100000000000247, 0.100000000000247,
  1.00000000000256, 0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255, 
    0.100000000000255, 0.100000000000255, 0.100000000000255,
  1.00000000000245, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244,
  1.00000000000254, 0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254, 
    0.100000000000254, 0.100000000000254, 0.100000000000254,
  1.00000000000268, 0.100000000000267, 0.100000000000267, 0.100000000000267, 
    0.100000000000267, 0.100000000000267, 0.100000000000267, 
    0.100000000000267, 0.100000000000267, 0.100000000000267,
  1.0000000000025, 0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249, 
    0.100000000000249, 0.100000000000249, 0.100000000000249,
  1.00000000000259, 0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258, 
    0.100000000000258, 0.100000000000258, 0.100000000000258,
  1.00000000000262, 0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261, 
    0.100000000000261, 0.100000000000261, 0.100000000000261,
  1.00000000000244, 0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244, 
    0.100000000000244, 0.100000000000244, 0.100000000000244 ;

 source =
  0.984804932153792, 0.0936887747126932, 0.0883219308441532, 
    0.101653616628478, 0.104190304978306, 0.0960705739442178, 
    0.101865315371057, 0.0905168693909131, 0.101722125465156, 
    0.103715066764544,
  0.971633170873509, 0.107203070824388, 0.0889566701318175, 
    0.101932103622956, 0.100380488128944, 0.096425276663493, 
    0.105195539764819, 0.0987048115474703, 0.102075617356411, 
    0.105811607136729,
  0.997285544966622, 0.10224183731164, 0.090657706545708, 0.108568682805694, 
    0.0966676155102172, 0.0974171830479638, 0.100720937442365, 
    0.0971998569568996, 0.0940299154601776, 0.110423176805444,
  1.00274777529196, 0.103157166335232, 0.0908581133199418, 0.108399431226952, 
    0.101385548512985, 0.0943743477162078, 0.101094301589055, 
    0.0937374450758755, 0.100354789174271, 0.103051782785613,
  0.983554134941522, 0.104554652659907, 0.0810215182965505, 
    0.114013014834488, 0.0943622679382315, 0.104061494621912, 
    0.102935011528312, 0.098434847343881, 0.0964091849555182, 
    0.106439720786692,
  0.959182797350487, 0.103881212528647, 0.093284679139645, 0.104654437354025, 
    0.105914874886979, 0.0983370219483563, 0.10038220280511, 
    0.0927837593956009, 0.101039971974924, 0.0991798112455935,
  0.986761803357476, 0.0994902306843554, 0.0908721140245701, 
    0.103002730019636, 0.104502760888792, 0.0975707114724476, 
    0.0992919832669225, 0.09991859576741, 0.0967326994131539, 
    0.106771764667479,
  0.965527012714905, 0.104376212022643, 0.0925171979183799, 
    0.104673102089275, 0.0926649158675021, 0.0993401985542511, 
    0.0993485643163904, 0.0958162282616226, 0.104747201305417, 
    0.10055309699646,
  1.00291981752586, 0.0971574731064237, 0.103473595660289, 
    0.0974035576963598, 0.10510638971514, 0.0949188652729292, 
    0.112073862916721, 0.0915969485037603, 0.095144048226096, 
    0.105449926844843,
  0.981705958680608, 0.103378286925711, 0.0950016313879153, 
    0.102819652085883, 0.0884017911600609, 0.0980988841672734, 
    0.104994256132328, 0.0949991824721936, 0.10443724425041, 
    0.0979510332565886,
  1.00812199977071, 0.0969455631361548, 0.0935023624806609, 
    0.108994102464054, 0.0924639717911049, 0.105861349552784, 
    0.101334388036189, 0.0961564088362944, 0.0944759388988835, 
    0.103377219411539,
  0.966044385168358, 0.103873032405053, 0.0911820462605042, 
    0.106209621260407, 0.0919964036849984, 0.103298760197144, 
    0.100824621550576, 0.0932958032634515, 0.0995483258786514, 
    0.104088911212376,
  0.99843350043955, 0.101412090506585, 0.0936869496648804, 0.113175177344318, 
    0.0866817307376796, 0.1023636773279, 0.101446999834287, 
    0.0933847958184368, 0.094779209307338, 0.110308997402841,
  1.02112884185471, 0.105046862188454, 0.0961552360903474, 0.106754651648581, 
    0.0907675285590619, 0.104454033948632, 0.103102925197339, 
    0.100520967299338, 0.0973675542718805, 0.100775021081974,
  0.991844531863358, 0.0990567685162587, 0.0972756853309114, 
    0.104787572089186, 0.0942795186414992, 0.105301938857449, 
    0.100578085086758, 0.0937444987740309, 0.0998694313847141, 
    0.100369160353784,
  0.987699868403273, 0.0988430088985149, 0.0942990896479416, 
    0.113481300257617, 0.0951855859213743, 0.103652205980268, 
    0.0980589497825107, 0.0975860209842827, 0.102534739345159, 
    0.105208593874045,
  0.988366515226378, 0.1029077120681, 0.0916373814978098, 0.109092953456372, 
    0.0991223166599373, 0.0953821969892996, 0.0992175587510897, 
    0.0998215171319427, 0.101441850064641, 0.0995373614338709,
  0.980390258784341, 0.0972494959742135, 0.0926230837019461, 
    0.0991016667428123, 0.101685197760749, 0.0936494054905756, 
    0.100749112434432, 0.0926113917925436, 0.100976630226657, 0.10900646747985,
  0.961334592014879, 0.0970687823591072, 0.088615554381664, 
    0.106189217950481, 0.0978875310908573, 0.0949267950067488, 
    0.104918422943155, 0.0933403515959989, 0.100909406548621, 
    0.101631577644992,
  0.97493136870604, 0.100625563432395, 0.0869278019800923, 
    0.0996150510141541, 0.0928235008046434, 0.100923177875655, 
    0.103565848568565, 0.0936855024374008, 0.0996665853093987, 
    0.107303869065547,
  0.9837850305492, 0.102107932614535, 0.0914307518627983, 0.104013070635289, 
    0.102367757761823, 0.101197956179153, 0.0976171517080918, 
    0.0921642111154666, 0.0917361946178126, 0.1026301665191,
  0.995605001058927, 0.102053593066703, 0.0923191862325898, 0.10247059931293, 
    0.0944760964848103, 0.102507003791029, 0.104077505534801, 
    0.0942847399107387, 0.103749373558884, 0.104107729773089,
  0.969050677797737, 0.1034654201738, 0.0829171907974395, 0.108300027078878, 
    0.103203718576089, 0.0948360815807032, 0.102264190112112, 
    0.0940569494909429, 0.0995790216073176, 0.106703793765482,
  0.976440004181433, 0.102483465513315, 0.0917305531501918, 
    0.104506165295508, 0.0997204479485125, 0.102701704994283, 
    0.104290056588119, 0.0968999197788235, 0.0963927696314476, 
    0.103489832810579,
  0.992802016607471, 0.101204736406198, 0.092164929448394, 0.106970712278851, 
    0.102751856576375, 0.103750254571375, 0.101689751114852, 
    0.0942864173697786, 0.0981685751477897, 0.100032084369397,
  0.989177837884752, 0.099669097331927, 0.0878422983661803, 
    0.105272069896372, 0.0981290215425117, 0.101170876896258, 
    0.103590922193714, 0.0944687638738297, 0.10675050382149, 0.106907165360344,
  0.962413834016745, 0.10729900141312, 0.0946627354388711, 0.106355553861522, 
    0.103108714984753, 0.0988048858673399, 0.102582642943431, 
    0.097510391535864, 0.103505775305022, 0.10595224184668,
  1.02382378970841, 0.101607036752099, 0.0835388948875953, 0.108117075459758, 
    0.0947972133664361, 0.0934843450456953, 0.0985136032557542, 
    0.0985368621588338, 0.0966863027383783, 0.104693904248956,
  0.958417747329014, 0.103285960371261, 0.0932288281366545, 0.10825961798412, 
    0.0967735410847719, 0.0961948899010086, 0.104930925244041, 
    0.0948237505886674, 0.104688388676818, 0.104243744480304,
  0.987274953628549, 0.099683157368269, 0.0903565044202512, 
    0.100610356813772, 0.0991619925438851, 0.10259092894634, 
    0.100589435557328, 0.0936058958211823, 0.10320742279623, 0.102468765951399,
  0.977721692595322, 0.0993870073575797, 0.0929605506406524, 
    0.104885975359902, 0.0979196835116193, 0.0931635231598495, 
    0.108892477264412, 0.0927690228970304, 0.0925885250655776, 
    0.109167089237824,
  0.958476981818758, 0.104823164880887, 0.0869606439549717, 
    0.109152838505121, 0.1010938689835, 0.0924557117908339, 
    0.106371276865536, 0.0912083267315794, 0.101283630321061, 
    0.105501948225434,
  0.952515103550448, 0.100443142560785, 0.0895211386652038, 
    0.107394703376934, 0.0939807279767763, 0.100737991151585, 
    0.107672754169272, 0.089142842590615, 0.101049649029773, 0.106479770143782,
  0.942047017264328, 0.105083147786066, 0.0847502061201557, 
    0.108737754775251, 0.0962602669796044, 0.102335173924305, 
    0.101485485542001, 0.099096256425536, 0.0985421155173633, 
    0.106838010895187,
  0.971886424054711, 0.103697526639773, 0.082450217694664, 0.108198052866541, 
    0.0981752210438431, 0.104651420059573, 0.0986816188316142, 
    0.0949166772205174, 0.0978824719716058, 0.107150479142247,
  0.975785772688849, 0.10838860718997, 0.0842744613623622, 0.111348830208919, 
    0.0964308160630643, 0.10320412007995, 0.102317096952037, 
    0.0964595724682114, 0.0974029452686923, 0.109291176734725,
  1.00005943567108, 0.0977131914208301, 0.0918623226556029, 
    0.104179675894552, 0.0935022943135018, 0.10243894203406, 
    0.101070213724587, 0.0947042617436466, 0.101631055242058, 0.10725427221926,
  0.99566769749999, 0.105061201916623, 0.0905524789973848, 0.107364519746076, 
    0.0963469739268191, 0.0976057535207727, 0.0992174604797254, 
    0.096668937088106, 0.103482374721587, 0.107264745996177,
  0.984143608885611, 0.103514012550863, 0.0835876212226326, 
    0.106484617608607, 0.0957216896229539, 0.0990507060915342, 
    0.10238390934181, 0.0921815274237658, 0.103209733696484, 0.105755372124323,
  0.987197849952706, 0.105479078673552, 0.0847412562095331, 
    0.103018864653518, 0.102580851209502, 0.0921235611467498, 
    0.107872619635858, 0.094142498419051, 0.0972008230520309, 
    0.105890506722023,
  1.00372726860624, 0.100492760518718, 0.0978395102431505, 0.10800045124667, 
    0.101486859078955, 0.0946419049455856, 0.107100144393301, 
    0.0925582197058649, 0.0983349740638723, 0.10862990769141,
  0.9933504934681, 0.101525528939811, 0.0803147848825951, 0.105308337347989, 
    0.0978082541465912, 0.104734599243612, 0.0974544337732925, 
    0.100655233358876, 0.10540962362947, 0.104896825231395,
  0.989956512707043, 0.0985792153142945, 0.0964773199352437, 
    0.103769161228533, 0.0991797781223381, 0.103972876652082, 
    0.0994467094822076, 0.0964767308502254, 0.100183604794487, 
    0.103482613090466,
  0.952688401861721, 0.096003414902295, 0.0993759914440725, 
    0.108769313908929, 0.0943037363624005, 0.106156178952991, 
    0.0996395794308675, 0.0954548996619614, 0.107769486114025, 
    0.0992241508037996,
  0.954053388318133, 0.100073807593975, 0.0936650475627276, 
    0.103635764240612, 0.0973140863977694, 0.102965563512914, 
    0.0999513560324575, 0.0973224824872635, 0.100918686029322, 
    0.104481719105407,
  1.00003703532259, 0.103078847074879, 0.0964228774534552, 0.106075151160225, 
    0.100087004521027, 0.0943188885120746, 0.105225741018952, 
    0.0926854935452743, 0.10733682077967, 0.100895673474479,
  1.0139734082295, 0.106676883612963, 0.0895945651190278, 0.108368283849029, 
    0.0959789621584264, 0.097795820104952, 0.102637465165047, 
    0.0981797317323539, 0.0940513660493444, 0.104230398191061,
  0.996731005809707, 0.0923977569576482, 0.09767443242001, 
    0.0987306077534504, 0.0987814850304212, 0.0991881938603743, 
    0.103889831264535, 0.0915470605156634, 0.0990321251843155, 
    0.100105682668005,
  0.940025005026449, 0.100841720635674, 0.0908869177848884, 
    0.106410201568832, 0.0983132069118878, 0.0995589534049027, 
    0.102162928288071, 0.0902717209716395, 0.0982159624157048, 
    0.104395885668104,
  0.975895358885207, 0.100718689419699, 0.0882503377224353, 
    0.107595464201988, 0.100237747898043, 0.0981999659578089, 
    0.0984376459312243, 0.095664883329551, 0.0987045058117938, 
    0.108384127564674,
  0.973153212801283, 0.107185283041656, 0.0860564463521476, 
    0.103864725746361, 0.0999965372883911, 0.0980114689408247, 
    0.104061936877114, 0.10000408220296, 0.101022700543951, 0.10730495632925,
  1.00464126880326, 0.10046441876185, 0.0895135992953225, 0.105527947749183, 
    0.0932285794005683, 0.0987557718610077, 0.0972299501919319, 
    0.0940039844674166, 0.0984255741535271, 0.104227782560423,
  0.992872180669526, 0.0998951062916611, 0.0888226175007147, 
    0.108877046221783, 0.0904517926259338, 0.107880245162758, 
    0.0986152596944393, 0.0980053868791762, 0.0968751482017902, 
    0.107196421850949,
  1.01134494080746, 0.0975879080445179, 0.0816962789297489, 
    0.106194389051193, 0.0955845419578689, 0.0998069525490813, 
    0.0953458001512099, 0.101504724877471, 0.0964603459641843, 
    0.104991130342522,
  1.02878757184882, 0.0989820015553989, 0.0930220442883803, 
    0.113074958878913, 0.0957634478240062, 0.102288946399385, 
    0.0994578599481901, 0.0944739960064242, 0.0966409558534755, 
    0.102075684769551,
  0.976847671886528, 0.108294039913032, 0.0869044622300634, 
    0.103759398494799, 0.0996559170603587, 0.10019718031071, 
    0.109015634051287, 0.0949601823570182, 0.0977206116122246, 
    0.107546665978352,
  0.958538992117635, 0.0993939921071114, 0.0871421739705726, 
    0.109559739014222, 0.0901439662152389, 0.103608620327415, 
    0.0971206935734406, 0.0983782329199913, 0.0922518129209291, 
    0.108208020440722,
  0.981872210834186, 0.099811417879141, 0.0896389702400007, 
    0.104738609406774, 0.0918764243609397, 0.101601238300503, 
    0.109004821432393, 0.0973920477285811, 0.0991720742846354, 
    0.106119625853548,
  0.965416928312579, 0.103242315418877, 0.097091608019919, 0.104439186159436, 
    0.0997090393203459, 0.102548591650005, 0.103563122026757, 
    0.0984678542515886, 0.103386146357247, 0.100935051649463,
  0.977914296291773, 0.102342054766937, 0.0911523976682517, 
    0.105163189267437, 0.0952246833200357, 0.0995065483877931, 
    0.10087777806624, 0.0967981816645242, 0.101625668531139, 0.101957711047463,
  0.991328497574221, 0.101869184864992, 0.0954776574157061, 
    0.104124178087385, 0.101880853167572, 0.101481161209597, 
    0.101316412157264, 0.0905568745387825, 0.0996422089491026, 
    0.099637526611431,
  1.00910825791638, 0.101488056954889, 0.0877262031488103, 0.111735674277099, 
    0.106124209548284, 0.0985706185442272, 0.101545279566808, 
    0.0926659583567155, 0.104275642123766, 0.100005761723418,
  0.976895786536091, 0.0990641522509226, 0.081991031988165, 
    0.107476025705598, 0.0993984739766507, 0.0967819840284943, 
    0.10605526656395, 0.0935565025083736, 0.102771934182828, 
    0.0976150387646272,
  1.00051076861208, 0.102479717992368, 0.0887591227059453, 0.101491842831803, 
    0.103093894809335, 0.104102016613495, 0.0994682349511002, 
    0.0980476896131505, 0.0972879455937195, 0.103223023657511,
  1.00453368670404, 0.0984532886448838, 0.089029123427684, 0.110776459535597, 
    0.102215201078719, 0.0984061259877287, 0.101211493597669, 
    0.0934238785800573, 0.101886741859106, 0.106332376304568,
  0.97630486687135, 0.0989241090610241, 0.0975591792211546, 
    0.108465948067285, 0.0984125765735969, 0.0947610004437861, 
    0.104605488294455, 0.0965363136484581, 0.101583496936203, 
    0.102058156691427,
  0.993500918065278, 0.0996164832599548, 0.0940932165998387, 
    0.11029176206546, 0.103010945329083, 0.100252167402195, 
    0.107741062221331, 0.0925341781758358, 0.0994917930351758, 
    0.104796673355736,
  0.979608976693719, 0.104905612342934, 0.103023462041668, 0.109149521069079, 
    0.094413638763561, 0.107438531599638, 0.101193867788803, 
    0.0964865825470698, 0.0996236627910508, 0.105706458967305,
  0.977415077218355, 0.0994580403268764, 0.0969035371399753, 
    0.0997688223769377, 0.108475009208907, 0.092768071689396, 
    0.104457025720031, 0.0964847039127858, 0.102040813257076, 
    0.106824503555519,
  1.00416321118563, 0.10124780007857, 0.0888844294998756, 0.110188024629638, 
    0.0984359748588474, 0.103247617900876, 0.101947352762093, 
    0.0960875902417675, 0.0999302938404655, 0.107339850938198,
  0.982022198662304, 0.103222555163672, 0.0807196062419703, 
    0.101621130713165, 0.0943890369257833, 0.0972350323126544, 
    0.103384023192336, 0.0987805467358254, 0.0957730541912857, 
    0.104755767233639,
  0.97760959307549, 0.0994641025491884, 0.0882903885504106, 
    0.107436394650298, 0.104165792470604, 0.0994631958539111, 
    0.106689215757643, 0.0913985787253077, 0.0987473920958107, 
    0.10421404090529,
  0.953233258238305, 0.099697952510334, 0.0890240871072824, 
    0.100850262459385, 0.101588834948596, 0.090874689685935, 
    0.102395644890792, 0.0941668972932187, 0.102079578174857, 
    0.103459160098125,
  0.986936667927081, 0.101651258336902, 0.0806396818091533, 
    0.110859374386735, 0.0884174856966876, 0.106920647194582, 
    0.100163343953398, 0.0951440136848801, 0.09646943000878, 0.103094523789385,
  0.973363898527197, 0.101835633972726, 0.090534327781806, 0.105984693307194, 
    0.103415135301368, 0.0913718591117477, 0.10636330458959, 
    0.0976034466338508, 0.0997956379931029, 0.105409810581965,
  0.955952302790603, 0.100212374940776, 0.095675183682529, 0.106170947754475, 
    0.101631734009234, 0.100870345656492, 0.103242914240582, 
    0.0974200845238418, 0.101002897972381, 0.103101063979264,
  0.985170870712743, 0.106969100619115, 0.0877669503749983, 
    0.104031493466296, 0.101161570182061, 0.100787085382036, 
    0.103580624333644, 0.0945296756953865, 0.0989871142575855, 
    0.102239902955088,
  0.97502523486209, 0.105754678097557, 0.0969424256685384, 
    0.0997037495158588, 0.0977281210154091, 0.101158421419312, 
    0.106534542422168, 0.0977989699154473, 0.0978861115484957, 
    0.101209160464682,
  0.962382399929706, 0.103832779301418, 0.10156942193105, 0.113334009584763, 
    0.096053704199541, 0.105124584375854, 0.0985113702226398, 
    0.0978808162968363, 0.102449117384034, 0.102868271682837,
  0.943543573643619, 0.100333566012261, 0.0923531836970572, 
    0.103210779680021, 0.104626861834925, 0.0922327786693389, 
    0.109929359890926, 0.0970332251798971, 0.0983839762563842, 
    0.107343785684853 ;

 source_phase =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wind =
  19.7834213155588, 21.3749369202483, 19.5048941243434, 20.9358862962633, 
    24.8535261361792, 23.5629878272439, 18.8111865682871, 20.9216450694202, 
    25.0509158970458, 19.0530470655968,
  26.1016035036898, 22.5795805483753, 21.9392735823064, 23.1974333593984, 
    25.4895391287202, 23.6334224908713, 21.7233244806447, 22.7119069485133, 
    23.3763982745132, 22.6412538367113,
  20.2804098594307, 24.1412623020681, 18.4885174708026, 19.6895185188231, 
    23.0795483602355, 20.4516202090494, 20.5180000376575, 23.7237028421857, 
    20.1474085863767, 18.9258416250284,
  20.8795132995587, 22.6328432090717, 20.4872915692096, 19.1896129994795, 
    24.3478856727997, 24.6380404602485, 25.0500374879553, 24.2204188152435, 
    23.6929834602246, 24.0293751550556,
  22.1973771921589, 18.6240665537242, 19.8510899886982, 21.0408278692619, 
    22.1817688729453, 25.3825759396857, 20.9599874586838, 21.3842942962745, 
    22.1768281183479, 20.513810204205,
  22.9510651118477, 19.6911002832542, 20.362754955908, 22.3591481370002, 
    26.2494607627871, 21.2187315000582, 20.9474660737749, 20.6290244963309, 
    21.5436264796061, 21.8714063445718,
  18.9519131881532, 20.3550077243242, 18.6931172774379, 19.6450630270883, 
    23.9904722931332, 27.0541994030575, 20.1651489627142, 20.3741833318033, 
    22.8901976959649, 20.7357877416816,
  20.7297190128901, 19.5560422895245, 21.3532825769671, 22.2760403245767, 
    21.6533625624899, 21.8496520149095, 20.5525138452258, 24.0189387252462, 
    22.5581084553832, 23.3683938046083,
  19.9485595539335, 23.0950782523567, 21.2005802182357, 22.7331469851878, 
    25.8052575592291, 25.7471163025467, 21.7924755139252, 21.8761583018766, 
    23.6556783801259, 22.7420846523912,
  18.7569906865681, 21.558266839881, 20.1735229304509, 19.9230378300906, 
    22.6282070851142, 25.3296284805052, 20.5367478562338, 20.3143640762417, 
    22.6841052195626, 21.5066812645182,
  22.690301070928, 22.8994970456699, 20.5884056464492, 19.7911245812188, 
    23.9042811813884, 23.7917299428444, 21.043603217831, 25.0231263853472, 
    22.7136415534366, 21.1751713440038,
  21.6151135554914, 20.2493459738598, 20.2564316221848, 20.2838339499383, 
    25.366077991826, 23.0597938412626, 19.3225757569434, 17.7906812108483, 
    22.1407302341943, 20.6585147380827,
  22.8685780351788, 23.2751735785102, 22.5956994587044, 21.1042291729448, 
    24.2385758613069, 23.9997289045794, 23.6764958382528, 25.5659786477662, 
    23.4899260686382, 21.1015239903733,
  23.7703589691923, 19.5182784700778, 19.7828947911803, 22.6036195304497, 
    27.5899913807006, 25.6574869540203, 21.6730534295881, 19.3052223670234, 
    19.9329743466101, 23.2451311177282,
  25.3792482326738, 21.604946470038, 21.8959529017763, 20.6170439602225, 
    28.3174089852057, 24.6239270723106, 21.8747920352692, 22.5759272067579, 
    22.6371709987449, 25.6693809138191,
  20.9600523705057, 21.0832521429001, 21.331474525387, 17.9377165245101, 
    25.019152505059, 20.9964784548614, 22.2396544769429, 21.3965468826336, 
    22.3266761773251, 21.8744677023707,
  23.2789466225271, 19.2180183115378, 17.7072771735491, 23.3640342820376, 
    22.7057218500969, 24.3358862982457, 23.1425229001992, 22.394099348731, 
    21.8852551701122, 23.7275800518554,
  19.2432499338955, 23.1207854907606, 21.810636828035, 19.1862499730884, 
    23.4348399565015, 22.6463385421307, 19.7502164712576, 21.2575355573656, 
    21.9369543518748, 21.6521967222628,
  23.0425163328272, 22.0317400703465, 24.0471290360478, 20.8678648153706, 
    24.9877648469608, 27.4582121380707, 24.0818081141521, 20.7915095179762, 
    21.7133397027969, 19.9369496810761,
  19.8897916338636, 20.3047385471954, 20.7276985643609, 21.3153976023967, 
    22.6748604021592, 22.5449618714206, 17.4451278762403, 19.6061648506022, 
    21.2633732652699, 21.4288249892872,
  22.6209318282509, 21.4874011685674, 18.789578751974, 19.4256189510477, 
    25.677213631235, 21.9916269999156, 21.804046310624, 22.1836173401298, 
    24.7054875481996, 21.1361331132115,
  17.5852453618893, 20.8096796760603, 20.8662831720319, 19.7290082516175, 
    25.5796319856725, 23.2318009197084, 23.1283042035846, 19.5120165365148, 
    22.5078636871479, 19.7972693735495,
  20.9072349842646, 23.6744836070178, 22.5454804243966, 20.0437366054498, 
    26.8400193758684, 24.9730343753821, 20.5464380040837, 22.245385493235, 
    25.5835897424107, 21.5860974223635,
  23.1025255001931, 20.9540728400828, 18.1741648980244, 19.8923034793996, 
    20.95026274998, 24.8755439797148, 20.2756619133753, 19.6268840663604, 
    21.0071804129712, 19.9418815997339,
  22.9295633734729, 22.4524346938718, 20.9888044672248, 23.2920951822708, 
    23.7628908584684, 24.6705570716303, 21.2486070128892, 20.175802401428, 
    20.4608756168679, 20.2133258660592,
  23.2989413762759, 21.4288400503514, 20.8647196498064, 21.6381780735322, 
    22.8228290771786, 24.0508640556587, 19.3658476292823, 20.5857992045396, 
    21.3743794280151, 20.9431463097047,
  21.5600110638292, 18.7600964227991, 18.935125837615, 20.636877436615, 
    23.2749456379626, 21.3823908871318, 19.7561195803346, 19.2018936274559, 
    21.4161995345083, 20.3502053814217,
  23.7498073175359, 22.998412532216, 21.2365785832895, 19.8419709286041, 
    27.6209528485147, 23.2202634373799, 20.9809058433692, 20.3819311903897, 
    23.160485801174, 24.8570109054371,
  18.984246648009, 20.6717962714018, 17.8284083170545, 22.6260864117023, 
    25.8255603505222, 26.4970244247111, 20.1118932190373, 21.8755416443022, 
    19.0353981591966, 18.7759270208256,
  20.0684107295973, 20.1515824706417, 19.3620336235171, 21.8590165070319, 
    24.4232322243951, 25.4967469953076, 22.0263209383708, 25.8654623634639, 
    25.0217677715524, 21.5795932905533,
  20.8620669700771, 19.8722522141707, 19.916492843869, 20.4395431124075, 
    22.2916649178225, 23.5590385839191, 23.0737488140098, 21.522931145102, 
    24.8008579172602, 24.5015839843473,
  25.4685115045088, 23.4547004028249, 21.542152553398, 21.8265461376617, 
    25.8679351342454, 25.2851890475787, 24.4129722573228, 23.5769476203696, 
    20.5497847158183, 25.6709254927266,
  21.561517689797, 18.0226503493777, 18.3378384668407, 19.3041650097476, 
    23.9464449800604, 22.9932505830307, 18.375405075196, 23.4637379686236, 
    23.2417803379612, 23.1411457704517,
  22.0283793464569, 22.1893249745422, 18.6604184293979, 22.1393560607841, 
    25.1216462637718, 23.462260772133, 20.5540805600772, 22.1907911068866, 
    20.0000286295402, 20.1776145766506,
  19.7841442865446, 19.4015433520828, 20.0025803552983, 19.2073475830857, 
    21.9170660590576, 24.3210995475758, 20.5419062749752, 19.1166688847929, 
    19.3062830446939, 20.2001926980517,
  23.8592831182352, 21.2948898697285, 20.2542012056384, 21.4915701269954, 
    22.5593513197812, 22.8897587677121, 21.8592399469025, 20.7735955378008, 
    22.7326290037784, 23.4002619189947,
  20.6662230039404, 20.7667802473159, 21.2564595349265, 22.9922259345168, 
    24.3917971146425, 24.2733377184249, 22.0441665102849, 19.531259774634, 
    20.8365152410248, 17.2787140447892,
  22.0216252411277, 24.1652259504095, 20.32431873512, 17.9833189391872, 
    25.1720757682342, 25.0550642985092, 20.9027771106528, 22.2295198928005, 
    24.1449721625632, 21.1229752086291,
  20.4536022010014, 20.3695317838347, 22.2465272640448, 22.8267799762675, 
    23.4463127576084, 23.4132784752047, 23.796780132773, 21.6847784280038, 
    20.0668250110103, 22.9674675510337,
  21.8208292178393, 21.0945616472626, 20.6629669412393, 23.4153991342513, 
    23.191481935867, 23.7320467665851, 19.780652238049, 22.1985537145181, 
    20.2936157243301, 23.2164233955687,
  21.8066934403246, 23.3089340149281, 23.3151085733394, 21.7535367031472, 
    23.8597001046467, 23.2872490324705, 20.8139802136552, 20.5799688692387, 
    21.0240018554822, 20.980942095243,
  21.4873885709527, 21.2993029477979, 22.1446184402709, 19.0689737961443, 
    24.1906921528617, 24.0465753940467, 21.5710722215052, 22.2949315775687, 
    21.0206968395772, 18.4188197341674,
  20.9643447121445, 23.2976398139152, 20.0578272393996, 19.8325657123015, 
    24.3265483669918, 25.5310240349818, 18.9670565786236, 20.1008615706072, 
    20.2197307017624, 20.8613882741379,
  21.2645629791237, 19.1268828776677, 20.4342131454917, 18.2609274566735, 
    20.66532440741, 24.0874292018476, 18.2358541427905, 23.8843743107101, 
    20.7265865985119, 20.3478788762404,
  22.0363200470396, 22.2811696193403, 20.4942866296828, 22.4223959460931, 
    22.2590282278384, 26.6191943327099, 22.7837747441078, 23.3931498053172, 
    19.6423475922688, 22.3041589453772,
  22.3606411113544, 18.3989590199739, 19.4131118322032, 23.4924172866558, 
    22.2961510536135, 24.2751967988868, 18.8940025028725, 22.4641460849638, 
    24.9615142907961, 23.3675186568998,
  23.6926921152653, 19.3441537776527, 20.8300399333158, 17.5674098277051, 
    23.1338215556784, 18.7770213714526, 18.298924936298, 21.452524283547, 
    20.6310079438982, 19.5488970210123,
  20.8318113919199, 21.1737348507528, 21.1418431605528, 20.8917857430678, 
    22.6501136381528, 26.6949376551286, 22.4146207396971, 20.7454080862955, 
    20.4879622441286, 20.5248968821201,
  22.1525014390339, 21.2122635753058, 18.5717192779706, 18.0653864533112, 
    23.693870810567, 22.6740942986071, 19.4471876520202, 23.7349365255431, 
    24.5573157615619, 22.9332344652366,
  21.5890830874341, 20.0794006009099, 20.8680149619297, 21.4182403058547, 
    23.3815199450305, 21.3193133590889, 18.966573935365, 18.6276918466402, 
    23.0519471841414, 22.4296784510591,
  23.0939179166903, 22.3257862121134, 19.5869684168222, 19.2331788712125, 
    25.3655196513867, 28.2710625333642, 22.9291443465534, 24.5993684241383, 
    21.5770880673461, 22.8210682811343,
  23.9168856535746, 22.0637540135255, 20.0297871393649, 21.1856580994117, 
    23.5170228604425, 22.5590344590885, 25.4484788666527, 23.8621199624062, 
    22.91144177778, 21.8382505573778,
  20.018003522442, 20.9875540400905, 19.935269846701, 18.8970838031295, 
    22.0480242132869, 21.7702775516866, 24.3695672569183, 19.902085652196, 
    23.0148247589002, 21.7033841324229,
  22.3008123215189, 23.2614210134525, 18.7377162571028, 20.8526606161724, 
    25.2978763662595, 25.0587528934217, 20.1960788220036, 17.535874931454, 
    23.0592142669411, 24.4059701008915,
  21.4389750257788, 18.0455509366148, 18.7005596167054, 21.5833640777449, 
    21.0893976739187, 22.5147777121078, 19.1605378881857, 23.4662598720356, 
    21.4470032345445, 21.2624735374525,
  17.4285252653796, 21.2574427567777, 19.6215306841312, 18.9922329061412, 
    22.8606984479898, 21.0651374005707, 17.985175322873, 21.0283880293816, 
    21.8149599448189, 17.9359000365268,
  23.3963890696894, 19.9817990877432, 19.307449165133, 20.7838457719383, 
    22.9529856076176, 24.0708616760719, 21.4800926386291, 20.5751990071104, 
    21.9134068388621, 25.3592220293074,
  21.3972617765864, 22.0962690573456, 21.8869113319922, 17.7675719024735, 
    27.2552976082639, 24.2939400203942, 22.8144621267217, 19.2399752873848, 
    22.3532243751254, 21.9798304581736,
  23.3783469421237, 22.3031099435685, 23.0087618438885, 22.1442005079262, 
    21.5397197238462, 21.8125908190417, 23.253539851858, 23.4796631821732, 
    21.181257160445, 21.2359323671332,
  19.1179285940465, 19.6772303865373, 15.6828751892208, 18.9705124529093, 
    21.6962638340846, 24.4048419622249, 19.3910429353694, 20.528881739317, 
    19.660483427517, 19.3751700383586,
  21.5943391299075, 19.1444916087499, 19.6118125212537, 19.8166529733051, 
    21.9870029130034, 19.7268964873411, 18.2998579586466, 20.015321742627, 
    21.5067252659213, 21.0858453286793,
  18.0087505539117, 22.643454066324, 19.6217953417406, 22.4130477843079, 
    22.9960626479449, 19.9090643526726, 21.9821867629336, 23.3683984403846, 
    19.0801270106913, 21.5603444023271,
  22.3276264570763, 22.0818886337134, 20.8793625103783, 23.5470567013673, 
    26.2734176732389, 24.2653473790403, 22.6465890589762, 21.0660339625865, 
    24.6142176538891, 22.2537654298826,
  21.9082339306264, 24.356063695429, 21.6599159647991, 21.869371700074, 
    21.020003770118, 23.5694462864432, 22.395220495918, 21.0572697081788, 
    21.683918724982, 21.1325666774503,
  21.9766075043467, 22.2419551505409, 21.5944711477169, 24.0110138924186, 
    25.7740553454722, 20.6602648861129, 20.7143869155774, 20.9739765232057, 
    21.0879710055023, 22.9233860008541,
  21.8746862309412, 21.3458534071748, 18.1083505424598, 21.2197208630805, 
    23.9502049924376, 22.5347500665727, 19.8673419796543, 22.1925822759365, 
    20.7359753447514, 18.8164778509411,
  19.8539983943516, 18.5257121291825, 20.2999945589101, 18.5815584902969, 
    22.7052831988667, 23.2228639534171, 18.1036047846562, 20.4847910589899, 
    21.5490989108365, 22.0921493793447,
  23.9412875724917, 22.0365398899722, 21.4341662299747, 20.8428300250908, 
    28.5934174232317, 23.8160958860942, 21.8298829624818, 24.0079565077527, 
    19.9327784171935, 24.4507953804553,
  20.96828275652, 22.0738120539839, 19.7681427737848, 17.4866376972965, 
    26.0795850696666, 22.7758373645906, 20.8357592546018, 23.9665619157978, 
    21.8564012993349, 22.1500825886632,
  22.5016428248309, 23.3112959074962, 21.4399223198096, 20.1871207417672, 
    25.4651905578958, 23.6451420055819, 19.451230322599, 24.6591953221823, 
    23.6546005351944, 21.0355999710231,
  22.7620313228309, 21.9434442557126, 20.8194315314356, 20.8320855441554, 
    24.6538823368526, 25.5885833656949, 22.8993833053727, 23.6197170904816, 
    25.9258805811369, 20.9561504912293,
  21.0747244443462, 21.7076693718179, 20.4318292159128, 21.2949424295247, 
    23.1144673296935, 24.60508724058, 21.6477048580857, 19.6436725912771, 
    22.4558002938395, 23.0283751426939,
  22.6848719232468, 21.4036001947904, 19.9883662996324, 20.2906950664386, 
    25.52731506305, 23.9804404773285, 21.544819125151, 24.2856725081757, 
    23.6379939422468, 20.6831751268682,
  23.3212716415537, 20.729936965919, 20.3934522487212, 20.1366128778877, 
    24.5441490443466, 25.2606414228321, 19.5606894062579, 19.137340878793, 
    22.3709799016828, 23.4815992629583,
  18.5548078673983, 19.7944929757683, 20.1829556125776, 19.1614540037596, 
    23.471886004453, 23.5945459059418, 19.5144936731612, 18.3275827762699, 
    22.0022517457591, 19.2257521404975,
  21.0691572230944, 21.2056144394924, 19.0567827702369, 19.9956764732369, 
    23.3544069574615, 23.1323658516111, 23.1506519102205, 21.173452935793, 
    24.516547972254, 25.1971728372186,
  21.4904808570759, 21.1994869071561, 21.9249973847693, 22.6855247153064, 
    25.023405861029, 29.2568050474308, 23.3107144233393, 22.4275359350139, 
    22.5445125155086, 21.6031105363902,
  19.3271683655299, 21.5165284579422, 20.6082864413544, 19.2668817138423, 
    24.2833602819263, 24.3136931144943, 22.638225110908, 19.935848288066, 
    21.934228114356, 22.1269296499483,
  21.842051579425, 22.9905303896846, 22.3731311634407, 22.2279069781631, 
    26.8686539083844, 25.3241584532736, 21.7968300246297, 21.8155790157438, 
    24.2195228589258, 23.8456102317852,
  19.7090742322303, 20.819895176926, 22.4769705197236, 20.0717330879359, 
    26.9201176011127, 23.9312232889809, 22.1324118194782, 21.0832562982629, 
    22.0226765562153, 22.0083792722252 ;

 concentration_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mean_source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_phase_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wind_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 concentration_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 mean_source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_phase_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 wind_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 location = 0, 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9 ;

 time = 41.666666666666667 ;

 advance_to_time = 41.666666666666667 ;
}
