netcdf wrf_bamex_00Z {
dimensions:
	Times = 37 ;
	x = 3 ;
	y = 3 ;
	x_stag = 4 ;
	y_stag = 4 ;
	z_amsl = 34 ;
	z_amsl_stag = 35 ;
	soil_levels = 4 ;
	ext_scalar = 1 ;
	record = UNLIMITED ; // (72 currently)
variables:
	int inityear(record, Times) ;
	int initmonth(record, Times) ;
	int initday(record, Times) ;
	int inithour(record, Times) ;
	float Z(record, Times, z_amsl_stag, y, x) ;
		Z:_FillValue = -999.f ;
		Z:description = "height AMSL" ;
		Z:units = "m" ;
	float T(record, Times, z_amsl, y, x) ;
		T:_FillValue = -999.f ;
		T:description = "Potential temperature" ;
		T:units = "K" ;
	float Q(record, Times, z_amsl, y, x) ;
		Q:_FillValue = -999.f ;
		Q:description = "Water vapor mixing ratio" ;
		Q:units = "kg/kg" ;
	float P(record, Times, z_amsl, y, x) ;
		P:_FillValue = -999.f ;
		P:description = "Pressure" ;
		P:units = "hPa" ;
	float U(record, Times, z_amsl, y, x_stag) ;
		U:_FillValue = -999.f ;
		U:description = "X-direction wind component" ;
		U:units = "m/s" ;
	float V(record, Times, z_amsl, y_stag, x) ;
		V:_FillValue = -999.f ;
		V:description = "Y-direction wind component" ;
		V:units = "m/s" ;
	float PRECIP(record, Times, y, x) ;
		PRECIP:_FillValue = -999.f ;
		PRECIP:description = "Run-time accumulated precip" ;
		PRECIP:units = "m" ;
	float MU(record, Times, y, x) ;
		MU:_FillValue = -999.f ;
		MU:description = "Total column mass" ;
		MU:units = "Pa" ;
	float MUB(record, Times, y, x) ;
		MUB:_FillValue = -999.f ;
		MUB:description = "Background column mass" ;
		MUB:units = "Pa" ;
	float MU0(record, Times, y, x) ;
		MU0:_FillValue = -999.f ;
		MU0:description = "Initial total column mass" ;
		MU0:units = "Pa" ;
	float ZNU(record, Times, z_amsl) ;
		ZNU:_FillValue = -999.f ;
		ZNU:description = "Eta values on momentum levels" ;
		ZNU:units = "" ;
	float ZNW(record, Times, z_amsl_stag) ;
		ZNW:_FillValue = -999.f ;
		ZNW:description = "Eta values on height (half) levels" ;
		ZNW:units = "" ;
	float P_TOP(record, Times, ext_scalar) ;
		P_TOP:_FillValue = -999.f ;
		P_TOP:description = "Pressure at the model top" ;
		P_TOP:units = "Pa" ;
	float MAPFAC_M(record, Times, y, x) ;
		MAPFAC_M:_FillValue = -999.f ;
		MAPFAC_M:description = "Map factor at mass points" ;
		MAPFAC_M:units = "" ;
	float T2(record, Times, y, x) ;
		T2:_FillValue = -999.f ;
		T2:description = "2-m temperature" ;
		T2:units = "K" ;
	float Q2(record, Times, y, x) ;
		Q2:_FillValue = -999.f ;
		Q2:description = "2-m mixing ratio" ;
		Q2:units = "kg/kg" ;
	float U10(record, Times, y, x) ;
		U10:_FillValue = -999.f ;
		U10:description = "10-m X-wind" ;
		U10:units = "m/s" ;
	float V10(record, Times, y, x) ;
		V10:_FillValue = -999.f ;
		V10:description = "10-m Y-wind" ;
		V10:units = "m/s" ;
	float TSK(record, Times, y, x) ;
		TSK:_FillValue = -999.f ;
		TSK:description = "Skin temperature" ;
		TSK:units = "K" ;
	float GLW(record, Times, y, x) ;
		GLW:_FillValue = -999.f ;
		GLW:description = "Downward longwave radiation" ;
		GLW:units = "W/m2" ;
	float GSW(record, Times, y, x) ;
		GSW:_FillValue = -999.f ;
		GSW:description = "Downward shortwave radiation" ;
		GSW:units = "W/m2" ;
	float TMN(record, Times, y, x) ;
		TMN:_FillValue = -999.f ;
		TMN:description = "SST" ;
		TMN:units = "K" ;
	float HFX(record, Times, y, x) ;
		HFX:_FillValue = -999.f ;
		HFX:description = "Upward heat flux at surface" ;
		HFX:units = "W/m2" ;
	float QFX(record, Times, y, x) ;
		QFX:_FillValue = -999.f ;
		QFX:description = "Upward moisture flux at surface" ;
		QFX:units = "kg/m2/s" ;
	float QSFC(record, Times, y, x) ;
		QSFC:_FillValue = -999.f ;
		QSFC:description = "Mixing ratio at the surface" ;
		QSFC:units = "kg/kg" ;
	float VEGFRA(record, Times, y, x) ;
		VEGFRA:_FillValue = -999.f ;
		VEGFRA:description = "Vegetation fraction" ;
		VEGFRA:units = "%" ;
	float ISLTYP(record, Times, y, x) ;
		ISLTYP:_FillValue = -999.f ;
		ISLTYP:description = "USGS soil type" ;
		ISLTYP:units = "category" ;
	float IVGTYP(record, Times, y, x) ;
		IVGTYP:_FillValue = -999.f ;
		IVGTYP:description = "USGS vegetation type" ;
		IVGTYP:units = "category" ;
	float LU_INDEX(record, Times, y, x) ;
		LU_INDEX:_FillValue = -999.f ;
		LU_INDEX:description = "USGS land use category" ;
		LU_INDEX:units = "category" ;
	float TSLB(record, Times, soil_levels, y, x) ;
		TSLB:_FillValue = -999.f ;
		TSLB:description = "Soil temperature" ;
		TSLB:units = "K" ;
	float SMOIS(record, Times, soil_levels, y, x) ;
		SMOIS:_FillValue = -999.f ;
		SMOIS:description = "Soil moisture" ;
		SMOIS:units = "kg/kg" ;
	float lats(record, Times, y, x) ;
	float lons(record, Times, y, x) ;
	float terrain(record, Times, y, x) ;
		terrain:_FillValue = -999.f ;
		terrain:description = "Land surface elevation" ;
		terrain:units = "m" ;

// global attributes:
		:times = "1-hourly" ;
		:contents = "profiles from WRF 4KM BAMEX run" ;
		:creation_date = "Thu Apr 27 12:38:54 MDT 2006" ;
		:TITLE = " OUTPUT FROM WRF V1.3 MODEL" ;
		:START_DATE = "2003-05-03_00:00:00" ;
		:WEST-EAST_GRID_DIMENSION = 501 ;
		:SOUTH-NORTH_GRID_DIMENSION = 501 ;
		:BOTTOM-TOP_GRID_DIMENSION = 34 ;
		:DYN_OPT = 2 ;
		:DIFF_OPT = 1 ;
		:KM_OPT = 4 ;
		:DAMP_OPT = 0 ;
		:KHDIF = 0.f ;
		:KVDIF = 0.f ;
		:MP_PHYSICS = 2 ;
		:RA_LW_PHYSICS = 1 ;
		:RA_SW_PHYSICS = 1 ;
		:BL_SFCLAY_PHYSICS = 1 ;
		:BL_SURFACE_PHYSICS = 2 ;
		:BL_PBL_PHYSICS = 1 ;
		:CU_PHYSICS = 0 ;
		:WEST-EAST_PATCH_START_UNSTAG = 377 ;
		:WEST-EAST_PATCH_END_UNSTAG = 500 ;
		:WEST-EAST_PATCH_START_STAG = 377 ;
		:WEST-EAST_PATCH_END_STAG = 501 ;
		:SOUTH-NORTH_PATCH_START_UNSTAG = 485 ;
		:SOUTH-NORTH_PATCH_END_UNSTAG = 500 ;
		:SOUTH-NORTH_PATCH_START_STAG = 485 ;
		:SOUTH-NORTH_PATCH_END_STAG = 501 ;
		:BOTTOM-TOP_PATCH_START_UNSTAG = 1 ;
		:BOTTOM-TOP_PATCH_END_UNSTAG = 34 ;
		:BOTTOM-TOP_PATCH_START_STAG = 1 ;
		:BOTTOM-TOP_PATCH_END_STAG = 35 ;
		:DX = 4000.f ;
		:DY = 4000.f ;
		:DT = 24.f ;
		:CEN_LAT = 40.00001f ;
		:CEN_LON = -95.f ;
		:TRUELAT1 = 30.f ;
		:TRUELAT2 = 45.f ;
		:GMT = 0.f ;
		:JULYR = 2003 ;
		:JULDAY = 123 ;
		:ISWATER = 16 ;
		:MAP_PROJ = 1 ;
		:MMINLU = "USGS" ;
		:SW_LON = -105.4442f ;
		:SW_LAT = 30.46228f ;
		:operation = "Conversion from old WRF input structure" ;
}
