netcdf perfect_input {
dimensions:
	member = 1 ;
	metadatalength = 32 ;
	TmpI = 60 ;
	TmpJ = 30 ;
	VelI = 60 ;
	VelJ = 29 ;
	lev = 5 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double TmpI(TmpI) ;
		TmpI:long_name = "longitude" ;
		TmpI:cartesian_axis = "X" ;
		TmpI:units = "degrees_east" ;
		TmpI:valid_range = 0., 360. ;

	double TmpJ(TmpJ) ;
		TmpJ:long_name = "latitude" ;
		TmpJ:cartesian_axis = "Y" ;
		TmpJ:units = "degrees_north" ;
		TmpJ:valid_range = -90., 90. ;

	double VelI(VelI) ;
		VelI:long_name = "longitude" ;
		VelI:cartesian_axis = "X" ;
		VelI:units = "degrees_east" ;
		VelI:valid_range = 0., 360.1 ;

	double VelJ(VelJ) ;
		VelJ:long_name = "latitude" ;
		VelJ:cartesian_axis = "Y" ;
		VelJ:units = "degrees_north" ;
		VelJ:valid_range = -90., 90. ;

	int lev(lev) ;
		lev:long_name = "level" ;
		lev:cartesian_axis = "Z" ;
		lev:units = "hPa" ;
		lev:positive = "down" ;

	double ps(time, member, TmpJ, TmpI) ;
		ps:long_name = "surface pressure" ;
		ps:units = "Pa" ;
		ps:units_long_name = "pascals" ;

	double t(time, member, lev, TmpJ, TmpI) ;
		t:long_name = "temperature" ;
		t:units = "degrees Kelvin" ;

	double u(time, member, lev, VelJ, VelI) ;
		u:long_name = "zonal wind component" ;
		u:units = "m/s" ;

	double v(time, member, lev, VelJ, VelI) ;
		v:long_name = "meridional wind component" ;
		v:units = "m/s" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
                time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		time:units = "days since 0000-01-01 00:00:00" ;

// global attributes:
		:title = "true state from control" ;
                :version = "$Id$" ;
		:model = "FMS_Bgrid" ;
		:history = "same values as in perfect_ics r1025 (circa Dec 2004)" ;
data:

 MemberMetadata =
  "true state" ;

 TmpI = 2.99999991876393, 8.9999997562918, 14.9999995938197, 
    20.9999994313475, 26.9999992688754, 32.9999991064033, 38.9999989439311, 
    44.999998781459, 50.9999986189869, 56.9999984565147, 62.9999982940426, 
    68.9999981315705, 74.9999979690983, 80.9999978066262, 86.9999976441541, 
    92.9999974816819, 98.9999973192098, 104.999997156738, 110.999996994266, 
    116.999996831793, 122.999996669321, 128.999996506849, 134.999996344377, 
    140.999996181905, 146.999996019433, 152.999995856961, 158.999995694488, 
    164.999995532016, 170.999995369544, 176.999995207072, 182.9999950446, 
    188.999994882128, 194.999994719656, 200.999994557184, 206.999994394711, 
    212.999994232239, 218.999994069767, 224.999993907295, 230.999993744823, 
    236.999993582351, 242.999993419879, 248.999993257406, 254.999993094934, 
    260.999992932462, 266.99999276999, 272.999992607518, 278.999992445046, 
    284.999992282574, 290.999992120102, 296.999991957629, 302.999991795157, 
    308.999991632685, 314.999991470213, 320.999991307741, 326.999991145269, 
    332.999990982797, 338.999990820324, 344.999990657852, 350.99999049538, 
    356.999990332908 ;

 TmpJ = -86.9999976441541, -80.9999978066262, -74.9999979690983, 
    -68.9999981315705, -62.9999982940426, -56.9999984565147, 
    -50.9999986189869, -44.999998781459, -38.9999989439311, 
    -32.9999991064033, -26.9999992688754, -20.9999994313475, 
    -14.9999995938197, -8.9999997562918, -2.99999991876393, 2.99999991876393, 
    8.9999997562918, 14.9999995938197, 20.9999994313475, 26.9999992688754, 
    32.9999991064033, 38.9999989439311, 44.999998781459, 50.9999986189869, 
    56.9999984565147, 62.9999982940426, 68.9999981315705, 74.9999979690983, 
    80.9999978066262, 86.9999976441541 ;

 VelI = 5.99999983752787, 11.9999996750557, 17.9999995125836, 
    23.9999993501115, 29.9999991876393, 35.9999990251672, 41.9999988626951, 
    47.9999987002229, 53.9999985377508, 59.9999983752787, 65.9999982128065, 
    71.9999980503344, 77.9999978878623, 83.9999977253901, 89.999997562918, 
    95.9999974004459, 101.999997237974, 107.999997075502, 113.999996913029, 
    119.999996750557, 125.999996588085, 131.999996425613, 137.999996263141, 
    143.999996100669, 149.999995938197, 155.999995775725, 161.999995613252, 
    167.99999545078, 173.999995288308, 179.999995125836, 185.999994963364, 
    191.999994800892, 197.99999463842, 203.999994475947, 209.999994313475, 
    215.999994151003, 221.999993988531, 227.999993826059, 233.999993663587, 
    239.999993501115, 245.999993338643, 251.99999317617, 257.999993013698, 
    263.999992851226, 269.999992688754, 275.999992526282, 281.99999236381, 
    287.999992201338, 293.999992038865, 299.999991876393, 305.999991713921, 
    311.999991551449, 317.999991388977, 323.999991226505, 329.999991064033, 
    335.999990901561, 341.999990739088, 347.999990576616, 353.999990414144, 
    359.999990251672 ;

 VelJ = -83.9999977253901, -77.9999978878623, -71.9999980503344, 
    -65.9999982128065, -59.9999983752787, -53.9999985377508, 
    -47.9999987002229, -41.9999988626951, -35.9999990251672, 
    -29.9999991876393, -23.9999993501115, -17.9999995125836, 
    -11.9999996750557, -5.99999983752787, 0, 5.99999983752787, 
    11.9999996750557, 17.9999995125836, 23.9999993501115, 29.9999991876393, 
    35.9999990251672, 41.9999988626951, 47.9999987002229, 53.9999985377508, 
    59.9999983752787, 65.9999982128065, 71.9999980503344, 77.9999978878623, 
    83.9999977253901 ;

 lev = 1, 2, 3, 4, 5 ;

 ps =
  101367.770704226, 101392.873808182, 101400.297346263, 101379.152078479, 
    101365.333810033, 101340.134757224, 101454.020680262, 101512.919261921, 
    101531.186212272, 101555.501346128, 101590.469709304, 101648.728566839, 
    101678.263488728, 101747.635060458, 101744.611322382, 101739.522170655, 
    101725.652785564, 101756.964709079, 101607.516378057, 101538.123497149, 
    101486.963711213, 101532.324896858, 101514.867667904, 101495.620891229, 
    101482.565662401, 101445.077648906, 101415.479326335, 101451.136623407, 
    101503.981886107, 101423.451109673, 101536.964761851, 101675.153995957, 
    101698.542280569, 101649.226739193, 101636.905486109, 101599.685109744, 
    101604.915148887, 101564.21006025, 101583.935487927, 101538.289027204, 
    101506.228080665, 101510.316257558, 101523.001164415, 101508.122877679, 
    101538.208671218, 101552.290272383, 101561.114573516, 101572.866055573, 
    101601.177062584, 101621.444130082, 101590.698787896, 101580.284462674, 
    101534.722582618, 101504.838048286, 101482.666660956, 101419.527332846, 
    101419.753676578, 101399.086389365, 101420.521873754, 101386.375861375,
  99877.5915625471, 99887.6142647717, 99962.6929788689, 100126.284844691, 
    100331.618552172, 100583.152593188, 100698.652660568, 100867.108476677, 
    101104.495359839, 101375.276435848, 101608.776995197, 101764.777214152, 
    101873.376923866, 101885.032328159, 101903.655555504, 101854.635846068, 
    101843.795421648, 101762.27708144, 101852.603996139, 101858.00746344, 
    101890.99615661, 101889.285154675, 101903.719811648, 101839.152104261, 
    101808.107580804, 101846.962872567, 101888.490265546, 101848.810221258, 
    101726.346492577, 101748.151428306, 101610.842793283, 101415.696396686, 
    101320.114843298, 101261.741603615, 101123.597934622, 101022.204740339, 
    100913.696162881, 100872.533821857, 100776.605994398, 100785.336601092, 
    100832.152726273, 100884.903821932, 100908.041893861, 100940.5080945, 
    100945.365365875, 100994.753776819, 101034.032019374, 101025.918416353, 
    100964.408690386, 100883.829176821, 100821.137573913, 100709.103238437, 
    100607.716237815, 100474.612880478, 100340.066955554, 100247.20024621, 
    100117.140284563, 100023.866601574, 99910.7849558445, 99877.414483341,
  100835.259214551, 100947.286218349, 101211.594773955, 101473.166765349, 
    101605.476571968, 101509.602836941, 101570.76972666, 101666.925328909, 
    101788.116198661, 101830.477539943, 101643.235538248, 101493.683844924, 
    101489.509691322, 101596.990803235, 101597.127629698, 101629.202698947, 
    101691.991238154, 102067.027736036, 102647.660629551, 102370.922692492, 
    101758.442912687, 101903.908144706, 101934.401115116, 101867.798058971, 
    101796.715491723, 101759.389357299, 101721.681437044, 101656.695743524, 
    101616.495679856, 101391.05762708, 101270.430705083, 101262.826706189, 
    101183.965372967, 101044.805374907, 100936.740596122, 100764.691282692, 
    100601.252944134, 100488.498538822, 100468.7007297, 100438.84181289, 
    100530.803725953, 100793.94353016, 101197.626491889, 101557.094993164, 
    101716.712235471, 101681.795004255, 101659.158344751, 101545.92280599, 
    101333.444883149, 101167.260863864, 101041.718346875, 101002.434871343, 
    100975.815854279, 100911.179865067, 100874.102745444, 100836.170306059, 
    100708.110367557, 100590.132661715, 100709.561736171, 100810.507526712,
  101423.020816594, 101541.33093813, 101394.108099772, 101186.627644603, 
    101152.076192662, 101375.554783274, 101540.540454652, 101480.738307286, 
    101003.241612971, 100338.612740892, 100212.910973379, 100696.967943804, 
    101167.019337019, 101625.259249205, 101903.198620136, 102307.838032302, 
    102587.581810629, 101909.99718286, 101149.764765608, 100564.164316738, 
    100316.809582315, 100361.932136576, 100486.341678843, 100778.999928315, 
    100988.073047758, 101112.409138434, 101273.000582, 101231.02890878, 
    101105.387989724, 101343.174221151, 101557.116530701, 101800.074088998, 
    101898.88811393, 101807.586826347, 101557.246300763, 101296.962564876, 
    101143.67433178, 101301.070388543, 101101.10319471, 100837.33901725, 
    100919.687803021, 101168.974050008, 101418.927206954, 101814.40738208, 
    102103.568662956, 102040.898047186, 101696.680309249, 101422.80938385, 
    101457.910649576, 101622.165492347, 101504.269426461, 101226.982926782, 
    101117.579514495, 100982.644292534, 100877.095211117, 100941.835645119, 
    100914.954387259, 101190.727449162, 101225.772709351, 101217.197374495,
  101467.034746459, 101473.826909203, 101101.071692285, 100984.995691921, 
    101407.327170372, 101523.856094527, 101229.917077935, 100492.304847692, 
    99667.2983950736, 99153.867884642, 99333.096300558, 99934.7870376973, 
    100913.927992225, 101853.86423335, 102151.893839731, 102094.384220495, 
    101407.804982111, 100440.50117437, 100062.359150516, 100265.587832364, 
    100475.18219066, 100912.275319173, 101055.679660479, 101040.258080699, 
    101181.401461599, 101314.007746102, 100907.59850139, 100559.591732, 
    101329.897627283, 102401.251916102, 102437.223635003, 101762.144777559, 
    101518.027900436, 101609.256344936, 101689.928090296, 101738.126584974, 
    101782.668422211, 101354.860033698, 100889.704528648, 100776.579439609, 
    101167.872805293, 101697.870086112, 102038.604705433, 102183.381829349, 
    102140.300016432, 101773.456476312, 101464.726764876, 101377.903705093, 
    101089.237055063, 100419.052365798, 99795.2052650686, 99959.4842427573, 
    100710.663942395, 101061.714779381, 101090.760288957, 101406.852215967, 
    101500.73735967, 100967.626193189, 100772.869494827, 101065.850086946,
  101487.271881388, 101682.372207506, 101628.69688351, 101715.837501708, 
    101579.399243475, 101271.378867068, 100895.619694606, 100293.276595668, 
    98812.2043311992, 97900.7409402231, 98035.0696937559, 98446.7524902733, 
    99586.0487826511, 100926.157120814, 101470.087758735, 101060.642741816, 
    100424.075837066, 99702.6144844476, 99997.1256690368, 100189.498540351, 
    100410.464440998, 101059.113582781, 102003.416766007, 101975.169763262, 
    101738.020642739, 101392.161766785, 100805.927190253, 101410.61990134, 
    102050.460086187, 101352.037881005, 100774.076420379, 101066.018364613, 
    101309.839380164, 101366.987413484, 101559.467222198, 101673.649450461, 
    101271.398865161, 100753.524296209, 100839.834184725, 101254.829596914, 
    101518.911614201, 101804.618558861, 101908.507831775, 101765.76497561, 
    101485.044065275, 101169.050161822, 100978.532387261, 100922.249262696, 
    100729.364187423, 100242.952992765, 99992.7960749712, 100617.571793145, 
    101326.345221941, 101687.049894544, 101647.275566685, 101314.455201202, 
    100698.570370131, 100613.991055866, 101031.659504025, 101402.627450367,
  100340.764731062, 100790.467731638, 100916.645103099, 100686.287011718, 
    100545.125437595, 100309.286030752, 100224.131744351, 100223.052859278, 
    99416.649550934, 98150.4708235121, 97520.2159036318, 97701.2026395559, 
    98528.1325745905, 99700.2136056783, 101254.930154293, 100450.027687942, 
    99920.1986415391, 99422.969909359, 99396.8224930495, 98855.4599284358, 
    99210.7635115862, 100054.80885307, 101249.174148007, 101674.259781018, 
    101911.469276472, 101912.575708799, 101831.830350305, 101809.918838379, 
    101104.007929141, 100125.114508286, 100038.046057966, 100521.151510429, 
    101265.917050542, 101460.358062994, 101444.860066443, 101128.687854544, 
    100555.974996767, 100136.736708359, 100066.078615218, 100313.008832317, 
    100780.505453134, 101060.658688834, 101235.122881953, 101046.153764686, 
    100749.841327051, 100372.402593113, 100168.416123724, 100151.809398166, 
    100312.949861592, 100385.002238059, 99985.3780431322, 99613.2267932097, 
    100108.455064937, 101216.852899195, 101179.556611559, 100440.175796875, 
    99634.8398379875, 99139.0231992855, 99227.8806747141, 100058.956866152,
  98544.358712095, 98689.3006729833, 99821.9297421771, 100245.092427638, 
    100344.536018638, 100040.352731388, 99937.6679936613, 99941.6420248065, 
    99769.7567243565, 99382.9519919167, 98866.2502995704, 98412.3128627245, 
    99603.3783649791, 98887.7718179021, 99345.8962361674, 100664.342047243, 
    100306.407387639, 99666.4701300724, 98659.2046421223, 97384.5754343224, 
    97659.9663609977, 98257.4684448801, 99730.7946626075, 100919.98209935, 
    101512.650014817, 101734.252445932, 101573.133498997, 101173.010772101, 
    100395.088524898, 99626.187472787, 99110.4452905994, 99414.9156969562, 
    99876.3400122065, 100164.505288943, 100165.769790271, 100208.813447073, 
    100255.064882324, 100153.531304353, 100069.29504974, 99659.1316532129, 
    99259.1661896494, 99589.4670118692, 100033.064382411, 100069.891147726, 
    99706.9997438015, 99131.2841629575, 98657.1231388426, 98562.1697310118, 
    98967.5365533955, 99897.2687854337, 100088.983685999, 100080.649683144, 
    99244.1094510832, 99415.4946108996, 100663.591123326, 100506.255191086, 
    100253.394011326, 100008.731059477, 100166.9016153, 99541.2557874444,
  99247.1452473733, 99655.9600515793, 100070.433733007, 100293.80736375, 
    99892.7618533859, 99399.6408186051, 99236.3907608618, 99226.8250667619, 
    99885.692330679, 100161.497269305, 100074.787873961, 99429.9082077884, 
    99708.2144849524, 100200.614571049, 99062.9064073116, 98787.9249399993, 
    100269.365931708, 100046.938080189, 99768.9083432015, 99273.5264065592, 
    98734.6018449256, 98479.8160340377, 98550.3120682736, 99548.5606544767, 
    100698.154473849, 100617.173742747, 99945.5602256026, 99533.5821130607, 
    99192.0543930857, 99361.4865556983, 99927.8459132992, 99492.9777397161, 
    98531.7928758805, 97830.6948980213, 98263.680541608, 98660.5743886692, 
    99123.8302099845, 99844.9829212932, 100184.104260952, 100132.74869286, 
    99726.990961706, 99190.1437794987, 99228.5436078409, 99392.4623450017, 
    99207.6479265738, 98955.9414196087, 98516.5091292987, 98371.8734310751, 
    98094.2826140641, 98882.9050198033, 100042.878159987, 100368.814478774, 
    99787.0830531109, 98448.4082110199, 97666.6315279308, 99515.7612378115, 
    100278.741592675, 100597.488635562, 100546.943481897, 99737.4682083957,
  98757.5610452282, 99013.4459590817, 100231.618105613, 100460.035589315, 
    99680.5127646308, 99835.3975731127, 99739.0696751352, 99221.8558795646, 
    99896.2794342925, 99788.8226841528, 99608.961401389, 100335.799473393, 
    100728.687149682, 100632.750715658, 99411.000381676, 98679.2339105665, 
    99597.086499679, 100595.187481002, 100694.485566988, 99855.0467650708, 
    99878.8407633944, 100376.692664772, 100082.191185124, 99745.2376047833, 
    99868.4639565826, 100134.434606967, 98991.1746102543, 98190.6985801759, 
    98091.4411452895, 98335.9231695905, 99600.3615155614, 100705.580182707, 
    99424.3730164667, 98810.353502505, 99940.17427071, 99821.5458868227, 
    98774.1026115183, 99190.8102482416, 100111.840731987, 100149.496886584, 
    99364.7362949182, 98612.4426241654, 98664.4308874923, 99629.7526221356, 
    100423.080812528, 99899.7728410348, 98745.1579804606, 99654.6036437522, 
    100093.749006079, 99270.1538062323, 99571.023561175, 100208.127363065, 
    99662.6532379777, 98008.415058096, 98115.1472264368, 98572.5576540532, 
    100012.690672266, 100743.147146997, 100573.103044464, 99795.2146095568,
  99141.7185269778, 99499.2030504014, 100411.488341282, 100393.285929054, 
    99718.6523672414, 99523.4325705074, 99520.2891977127, 100043.036754688, 
    99561.1796001631, 99784.2961840806, 100647.697325543, 100304.768049332, 
    100257.945494726, 100117.05647296, 99469.9682885337, 99454.721295364, 
    99773.2380783231, 100629.787197797, 101050.315390249, 101015.214597674, 
    100077.52851354, 99331.9925412841, 99619.0137650654, 99894.4863969149, 
    100221.98960233, 100109.816667805, 99687.1407911986, 99273.4174754187, 
    99536.7120135074, 99698.2557688867, 99875.5264193326, 100161.135756606, 
    99923.3249420484, 99975.4936610296, 99651.8950222084, 99420.9390128133, 
    99373.8865119217, 99724.6805861866, 100103.638587844, 99926.4876403971, 
    99626.5160939094, 99278.8524667539, 99380.7815082192, 99867.8650738085, 
    100188.759738565, 99946.1978826811, 99940.0026808292, 100055.65602387, 
    99797.4875527851, 99362.1590907375, 99690.3148447659, 100010.668887052, 
    99637.0439075242, 98968.7049819795, 98843.7247594138, 99595.6188720583, 
    100064.855098556, 100596.712726853, 100303.675456712, 99595.3188294841,
  99586.6140749389, 99765.353597899, 100018.811155194, 100031.861385568, 
    99827.3680231332, 99837.4937686008, 99859.7111345472, 100166.22905581, 
    100426.432571108, 100358.274628034, 100049.521249384, 99768.4929409968, 
    99762.5147252348, 99823.8115389636, 99943.7949788439, 99933.2636884016, 
    100352.044333251, 100677.839703854, 100508.259445683, 100027.449548006, 
    99615.5029503261, 100156.87270349, 100360.429524604, 100396.700157162, 
    100490.669010808, 100366.361099778, 100089.989053854, 99194.5284091224, 
    99296.9547007793, 99982.6183065264, 100220.293929226, 100330.964998569, 
    100281.942569574, 99878.0808149725, 99402.2670416429, 99278.3741404382, 
    99580.0100756578, 99902.6809781266, 99973.4450625572, 99886.6411494151, 
    99622.4371667231, 99659.0693761259, 99871.1524341032, 100106.021302105, 
    100261.053031446, 100167.932229167, 99896.9050501769, 99671.3883211826, 
    99682.8864755984, 99904.1635460655, 100065.607784, 100085.664848502, 
    99844.5489656301, 99366.0049569347, 99294.1756941545, 99563.2411119076, 
    99974.7074504224, 100224.452501004, 99943.2493010716, 99609.3808039517,
  99426.6964675892, 99604.3900158976, 99779.5393928274, 99797.1183514588, 
    99854.3102224208, 99941.8440565793, 99930.4237795695, 100057.940837959, 
    100040.299031645, 99999.3677758834, 99843.3454102011, 99628.2326106627, 
    99790.2209364786, 99864.6221548251, 99928.8384467891, 99979.7027445749, 
    100099.853861441, 100179.77924154, 100040.951000174, 99718.3666058407, 
    99777.374932597, 100096.865282023, 100167.782086625, 100151.216291558, 
    100269.10872308, 100212.759155528, 99735.8320093587, 99617.6713579957, 
    99732.6726153271, 99802.9934690629, 99947.2715171596, 99972.8491964149, 
    99915.8150763411, 99645.5676028462, 99574.9790479441, 99579.6304532626, 
    99623.9794116632, 99688.5875365606, 99775.1065827092, 99736.7938718794, 
    99577.7216590761, 99581.5044784648, 99705.7046582978, 99871.6621463076, 
    99912.8995573269, 99852.9909664566, 99660.9790563568, 99648.4787204039, 
    99686.5644591461, 99747.689379526, 99823.0489390276, 99807.5412048921, 
    99505.1676323083, 99331.7865365176, 99522.9155751704, 99664.995850213, 
    99782.2831449803, 99849.8266622979, 99764.0157768092, 99522.9782667834,
  99475.9346824599, 99442.2537471799, 99624.7032129421, 99666.1638059553, 
    99732.3080070136, 99810.9596423081, 99874.6745361617, 99916.8611872471, 
    99905.3159815985, 99859.2967687821, 99514.1904487257, 99541.1993212169, 
    99619.6307693276, 99676.9051402843, 99734.7330275634, 99812.9224554937, 
    99846.5418802911, 99806.9470358266, 99570.4949107364, 99487.0150952651, 
    99603.1046104374, 99674.3832655801, 99877.8101738853, 99827.3279387119, 
    99861.5636504537, 99680.8190090478, 99507.0412763744, 99522.9499868861, 
    99579.0792982557, 99647.965290123, 99680.9566022676, 99663.4874275223, 
    99560.3124313442, 99488.8429508459, 99458.9023225243, 99482.942821791, 
    99484.5289239132, 99498.7478624408, 99551.3295085563, 99563.9563525733, 
    99485.9244520658, 99462.0546088966, 99534.4678708693, 99580.0319927614, 
    99594.1490088261, 99517.5446620687, 99488.9477141937, 99511.6203732378, 
    99588.7410952153, 99607.4211936666, 99599.1735041119, 99553.7074670975, 
    99424.0032822325, 99355.5367366527, 99414.8381176067, 99485.3399926638, 
    99553.1492110412, 99583.1218743384, 99542.0755619071, 99494.0195206507,
  99377.2342345128, 99460.3160325202, 99481.2471476489, 99565.7548778825, 
    99690.9355813785, 99617.6819427524, 99575.8476459296, 99599.6989692572, 
    99666.2029253385, 99576.6522994286, 99424.9664013635, 99425.3880153383, 
    99462.2724073902, 99503.3769943662, 99549.6039164156, 99536.1163749675, 
    99552.6842214088, 99533.5988075052, 99367.3165337234, 99413.37507826, 
    99487.620137601, 99508.3354507145, 99555.6325036488, 99483.9679729947, 
    99574.244927021, 99441.1376192773, 99403.5517617705, 99430.7237081249, 
    99467.3465258339, 99513.5257219166, 99523.3204116193, 99494.2468887858, 
    99399.2725863542, 99339.831633006, 99371.3709972565, 99365.7129190774, 
    99362.3302327681, 99367.3743121645, 99424.4449852528, 99443.6446992234, 
    99425.5501294415, 99404.2303473051, 99341.8613867884, 99373.1520950928, 
    99391.370641174, 99340.3934479816, 99351.2950625246, 99396.9353093454, 
    99382.738679273, 99370.500473743, 99422.2907425442, 99436.9646427041, 
    99360.2679065327, 99283.4286709923, 99340.3811553061, 99369.3676354894, 
    99373.0539914791, 99380.6950240985, 99373.4213694766, 99408.3285206879,
  99437.7682735797, 99399.120819699, 99431.8118061492, 99496.2047429543, 
    99524.3581499285, 99480.6114290912, 99431.7046685106, 99606.7079834506, 
    99726.1671660606, 99637.6157893017, 99458.9336649612, 99351.5527114311, 
    99383.0232858544, 99392.710032923, 99399.8396253563, 99456.5187346168, 
    99436.4985045669, 99413.8742428583, 99398.6172107663, 99392.4769195547, 
    99393.3094834952, 99464.5044503136, 99453.7464424903, 99395.75300824, 
    99362.6183631951, 99424.5382523857, 99468.0764324437, 99441.5199804969, 
    99523.202610338, 99556.458538864, 99553.6412032185, 99548.9026161279, 
    99455.2162918807, 99387.1497267861, 99348.1209383597, 99372.4407159746, 
    99353.6893286855, 99352.5214407236, 99332.8877469359, 99374.2565234476, 
    99410.7176816445, 99406.6843484317, 99339.7667257293, 99350.4440523598, 
    99386.5685458179, 99368.2595136435, 99348.520724666, 99337.8862010595, 
    99349.0221657919, 99330.4363081256, 99329.7262401636, 99353.0658281788, 
    99325.1968218866, 99318.4021020722, 99340.2043668121, 99362.6843090074, 
    99330.4609925397, 99317.4065489921, 99400.2558772329, 99395.9009856374,
  99666.0210475162, 99622.6422791418, 99432.2026685765, 99505.4081651772, 
    99533.0867187322, 99540.0438046382, 99606.5746624605, 99628.2618615124, 
    99631.0101137197, 99543.548980813, 99422.857118915, 99437.643570132, 
    99443.6745069505, 99457.6949804824, 99437.6403237358, 99387.5069680413, 
    99423.6240653238, 99477.4698826959, 99498.9481097385, 99496.9172755928, 
    99499.6340943334, 99511.707127889, 99521.4644354649, 99486.4366995652, 
    99477.631370301, 99511.9587474304, 99610.9806028831, 99713.5796628712, 
    99725.1808168977, 99794.8415389921, 99893.1286610094, 99793.7347022421, 
    99512.6138586529, 99430.7875554646, 99432.8489091837, 99428.3361197118, 
    99469.0658063434, 99495.6163339207, 99471.3187228663, 99546.4435653993, 
    99517.7369408857, 99497.5321638974, 99448.8926588494, 99465.9081094537, 
    99504.3693064707, 99517.856848781, 99478.9805544918, 99449.5802486286, 
    99392.0470288237, 99395.2805708837, 99363.7775525071, 99414.7170141319, 
    99458.2258013463, 99478.002486703, 99446.9792307183, 99440.8677061989, 
    99444.253293084, 99434.2944533562, 99440.8775750944, 99527.1679054834,
  99809.6174653381, 99925.8036512262, 99784.2595798815, 99710.8757740127, 
    99585.2611477978, 99661.3995853892, 99810.0431088806, 99968.034681222, 
    100108.764408175, 99923.9411863695, 99574.4733654081, 99479.4964694758, 
    99635.0060776168, 99618.6238348608, 99544.5420511328, 99478.9193170757, 
    99542.001163753, 99603.3093098728, 99628.8334784651, 99654.1764619156, 
    99649.3097375919, 99729.4995655691, 99692.7517889989, 99632.7934656084, 
    99530.139519836, 99627.5984806389, 99828.4966620661, 99933.4249444298, 
    100058.078879051, 100127.324386849, 100208.062703627, 100200.730259247, 
    99827.1095215737, 99664.3762636606, 99520.1830094318, 99647.7193015859, 
    99750.6429848038, 99820.4855284869, 99865.4667357053, 99782.5617780853, 
    99675.1056723947, 99581.9791383274, 99544.2846553966, 99642.8915374691, 
    99736.9370128966, 99752.2822649746, 99731.8202412755, 99640.2285136725, 
    99543.7840450757, 99488.3018650658, 99510.1241236242, 99571.720680558, 
    99685.7353093131, 99687.6290274006, 99730.2994560245, 99795.5785004052, 
    99723.9580188709, 99655.8093567763, 99526.3912744671, 99732.1071401083,
  100235.234751438, 100352.740963064, 100392.408737877, 100002.838668482, 
    99800.5624610546, 99967.9879902889, 100178.549828612, 100470.209254521, 
    100578.404220079, 100579.018117366, 99905.4448001358, 99553.1769813503, 
    99753.0674480867, 99843.7135003727, 99838.8304687138, 99874.0755701445, 
    99909.700664549, 99799.8387372419, 99817.2844471432, 99750.5572788267, 
    99854.2411474507, 100032.270090307, 100148.514301993, 99927.4619702057, 
    99765.2086517114, 99774.3411976468, 99918.0457371396, 100058.756839744, 
    100214.314745054, 100409.984879954, 100529.35078014, 100661.036165203, 
    100366.639611826, 99874.4036955332, 99591.5596259605, 99740.0909765203, 
    100000.108408571, 100084.887322291, 100234.167280145, 100199.32071004, 
    99901.4159597852, 99745.6588659569, 99721.7323016417, 99874.0424142854, 
    99996.8505946898, 100045.892287149, 100103.147212128, 100050.724374108, 
    99869.118258961, 99873.2214681371, 99918.8655864766, 99953.3397333738, 
    100012.319485338, 100087.922784237, 100186.416244241, 100227.558415343, 
    100211.151952845, 100004.64384107, 99770.2144949654, 99901.6473268897,
  99297.2430712424, 100453.108190212, 100914.713973571, 100690.982741905, 
    99534.556555409, 99481.1282077334, 100298.683333196, 100748.232452952, 
    100953.536010385, 100901.517832794, 100370.524224386, 99197.650787689, 
    99320.8890181214, 99790.9045421406, 100470.236904185, 100618.777972818, 
    100522.458042742, 99972.1105125899, 99585.3099332579, 99851.6294552012, 
    100287.521904821, 100685.762094011, 100811.177520234, 100475.848593019, 
    100070.533492772, 100181.497401456, 100002.073525002, 99595.171793963, 
    99438.3338297249, 99880.3640651751, 100355.573981937, 100684.242674012, 
    100750.646488144, 100268.726759628, 99687.900382786, 99570.6641274669, 
    99567.3458705284, 99516.709627077, 99836.0384915363, 100272.439201677, 
    100365.383208825, 100125.775827402, 99790.189021425, 99714.823391855, 
    99879.9058559077, 99984.1375635585, 100310.443639599, 100596.965724662, 
    100502.696828392, 100595.311772158, 100797.97257058, 100695.253135963, 
    99966.1595801758, 99773.3942464526, 99842.8915736947, 99985.8113932913, 
    99998.099216826, 99858.7318151201, 99769.9954925593, 99354.1798179167,
  99573.9722201084, 100681.147896589, 100348.863154685, 100489.518290498, 
    100413.059453473, 99956.8598394607, 100365.540429216, 100235.951938995, 
    100156.195005276, 100299.628864971, 99911.8563727018, 98908.4940874334, 
    98452.9036907228, 99801.0669751056, 100777.178219831, 100993.920899274, 
    100436.049996623, 100150.329689777, 99897.1221367672, 100034.37554229, 
    100665.526451471, 101320.455949324, 101578.298446478, 101033.485222529, 
    99987.3462485225, 100068.820109978, 100163.475728823, 99635.6809521345, 
    98766.7137583629, 99188.0771796296, 99951.3634879157, 100167.346097966, 
    100269.472043347, 100139.597498088, 99734.9912918693, 99155.3325053136, 
    99136.0079416192, 99948.6075566431, 100414.312754034, 99967.0832310889, 
    99837.2650161483, 100179.818504432, 99932.722892883, 99338.5540560109, 
    99757.0735514839, 100076.377089497, 99661.8945991761, 99824.2891152554, 
    100470.025218964, 100784.445797287, 101285.438692033, 101700.413089049, 
    100573.706893362, 99656.9680145644, 99778.7076901393, 99452.2085869628, 
    99670.9622876917, 99140.0118464022, 98057.4968316994, 97813.4380259641,
  100192.915489418, 100112.359583383, 99464.6335100216, 99029.1274661899, 
    99398.4835914899, 99257.5610540841, 98476.6942361604, 99244.8684635721, 
    100256.779222467, 99997.2425536565, 98924.780505567, 98200.6618252625, 
    98292.8751944048, 98915.7178365139, 99924.5605428307, 100744.78726113, 
    100365.423877892, 99000.9249787601, 98074.6739633839, 98631.7402543693, 
    99924.8883826207, 100868.022058439, 101281.902280753, 100995.945077368, 
    100058.542863222, 99123.888928719, 99583.1618437399, 99277.962309127, 
    99414.0826101821, 100106.199733058, 99797.1118081949, 99637.5656163773, 
    99447.5430990781, 98905.6857823088, 98042.8602253618, 98072.5029766223, 
    98901.9614487479, 99933.3063921524, 100519.335981928, 100089.913341084, 
    99725.9500481444, 99950.474284551, 99233.0628788342, 99213.0280775007, 
    99269.1754740383, 99933.0445441085, 100519.982899982, 100642.802384029, 
    100821.338280245, 100539.407148565, 100303.632622098, 100215.277933812, 
    99608.2433871036, 100517.585675269, 100493.486200501, 99488.0976513871, 
    100565.048619657, 100740.703705219, 100532.94888332, 99962.8892959854,
  99817.9204536574, 98203.8181683083, 97465.3556056229, 97339.4893124073, 
    97323.200866782, 97734.2909941952, 98912.0086866051, 100080.532381813, 
    99890.7638351601, 99216.0730135349, 98423.9444354446, 97948.4481589913, 
    98457.3628959782, 99239.1068655063, 99897.2238042469, 100904.857517357, 
    101298.775830648, 100428.99442328, 99490.3968317561, 99184.9062004047, 
    99457.5072029464, 100082.645213225, 100131.58671051, 98611.5692535348, 
    97873.8184088105, 98789.0796847017, 99164.8074245096, 99496.2123431385, 
    100425.133152176, 100235.240636285, 100100.099050058, 99618.6516406623, 
    98752.0881974538, 98420.3791648431, 98434.9498526523, 99050.2872925873, 
    99910.8022070395, 100515.804762386, 100629.177775052, 100581.438021223, 
    99965.418644846, 99664.2759917178, 98455.0241656553, 97935.6303647777, 
    99172.3529629006, 100729.647716642, 100977.54697589, 100904.144950452, 
    99887.4765059203, 98964.5227842923, 98670.0371393585, 98515.5790722415, 
    98297.7942261822, 98401.7060892034, 98652.9521728554, 99848.6345896842, 
    100644.050666305, 100672.985652925, 100842.850314112, 100400.82055617,
  99883.9053099441, 99530.9809561124, 99230.4656985357, 99314.2889015209, 
    99368.3398386086, 99916.9722738163, 100176.333475998, 99887.921637626, 
    99459.0294878041, 99421.2317583286, 99567.7837240583, 99666.573799878, 
    100096.968116381, 100528.316764561, 100901.747117302, 101189.711729895, 
    100855.837737586, 100569.087363485, 100378.535604926, 99917.4095558593, 
    99585.4513831501, 99142.9135335805, 98597.8525595012, 98537.922202911, 
    98822.9973725934, 99079.5119275085, 99503.1142513123, 100370.926062389, 
    101022.600756592, 100976.868787022, 100997.57401868, 100907.489973728, 
    100755.452277711, 100723.600885166, 100887.366099888, 101298.004779257, 
    101511.797533779, 101385.263014662, 100704.610281971, 100074.651323954, 
    99267.7606625547, 98240.4894934081, 98654.521191415, 99528.1399688416, 
    100635.906072192, 101199.317712804, 100988.054067601, 99742.1038832271, 
    97943.6076017368, 97915.0601978025, 98725.7943180399, 98341.8061136186, 
    98177.1542998989, 98599.9750840132, 99266.824917966, 100195.825107209, 
    100590.472718454, 101051.027839126, 101080.746284877, 100552.833133044,
  100163.860837013, 100403.266307328, 100713.617835821, 100825.87178445, 
    101054.832588777, 101108.15688574, 100886.992124653, 100440.652915284, 
    100003.462870854, 100150.714959724, 100631.360749325, 100837.487884535, 
    101063.335071593, 101304.243713027, 101266.268125635, 101049.687286855, 
    100471.739641161, 99869.94148046, 99729.2590546166, 99455.2444811708, 
    98978.8945590293, 99164.4677765886, 99404.0152329396, 99824.5959226034, 
    100129.951175871, 100448.305538078, 100790.770382578, 101072.738804203, 
    101052.981488212, 101025.35722208, 101017.323057891, 101225.502543652, 
    101477.314076041, 101766.530803912, 101955.990086773, 101992.278720863, 
    101835.364062914, 101081.245586394, 99914.6291914258, 99465.1954378913, 
    99475.9926015543, 99457.2334347865, 100361.517467516, 101162.371891165, 
    101369.722927918, 101301.507596342, 100855.52001779, 100039.250655291, 
    100384.609080218, 100509.93838921, 100210.858855374, 100197.080822573, 
    100262.253667785, 100253.641695029, 100306.207071299, 100632.566282371, 
    100700.973312791, 101118.675706203, 101300.254907602, 100689.145044051,
  100635.210907105, 100579.315391903, 100901.99143477, 101326.108296726, 
    101771.745514515, 102050.853973272, 101929.412451578, 101413.715896346, 
    100791.888017013, 100614.620147676, 100883.888582178, 101124.53219995, 
    101317.360248884, 101522.731919643, 101586.115588847, 101149.48256439, 
    100547.709399836, 100108.162231112, 99857.3646163274, 99927.7406770393, 
    100170.064750065, 100473.169054448, 100898.530090012, 101211.997491002, 
    101511.526345087, 101650.901706361, 101757.981311189, 101654.214612014, 
    101522.679911445, 101306.713728089, 101169.300537099, 101130.589723866, 
    101174.051470642, 101056.576079812, 100929.202990035, 101303.725211239, 
    101693.403333631, 100998.071179424, 99801.0804779928, 99322.6404619222, 
    99830.4499908118, 100619.698475525, 101417.349444881, 101839.510340657, 
    101759.496394784, 101753.587228238, 101652.000808441, 101246.401687246, 
    100656.235011365, 101070.022434988, 101419.140172405, 101520.295703402, 
    101308.180031585, 101063.294534538, 101069.798057623, 101093.397744324, 
    101071.508625457, 101096.676319389, 101109.992310772, 100917.089059955,
  101255.26681936, 101038.963845936, 101173.118457052, 101385.364519449, 
    101629.271571971, 101906.65699268, 102240.472343702, 102378.256505018, 
    102069.266737211, 101531.025975461, 101159.346058617, 101060.103132229, 
    101141.371903903, 101364.118804461, 101445.34474989, 101311.585241629, 
    100914.038728126, 100529.291254298, 100415.985195412, 100467.845978725, 
    100652.824920668, 100944.336922692, 101151.726011635, 101480.864923899, 
    101697.551219415, 101868.656639883, 101872.455423549, 101813.472654681, 
    101648.207927892, 101518.412132382, 101447.286500305, 101416.579428022, 
    101255.590494722, 100976.939110833, 100749.576567253, 100971.534901818, 
    101503.203680994, 102108.932381094, 101633.394692908, 100637.083297144, 
    100581.149238468, 100724.008506194, 101041.414663547, 101377.058007808, 
    101577.37015478, 101469.58455254, 101195.482682526, 101289.822614492, 
    101863.57242388, 101940.724664942, 101845.922180658, 101901.96360117, 
    101991.300763144, 102090.595070613, 102188.142254396, 102252.962389155, 
    102239.605456907, 102122.943992955, 101813.591539231, 101505.409193209,
  101595.305768745, 101340.443944703, 101180.720713194, 101131.562267007, 
    101229.614193742, 101458.39415883, 101689.975775873, 101920.94893637, 
    102076.371890314, 102051.231635174, 101739.704441462, 101330.393720308, 
    101103.80485368, 100992.038054694, 101022.110688267, 101142.670851895, 
    101301.737432109, 101227.170079838, 101069.433450872, 101001.671861582, 
    101058.908153677, 101114.851956788, 101228.374350457, 101321.196714753, 
    101453.138295347, 101437.669319627, 101283.339663319, 101112.348726689, 
    100975.451958459, 100786.073742566, 100745.738749091, 100807.268186341, 
    100932.860493195, 101069.067540188, 101176.886761295, 101317.767121215, 
    101487.25212048, 101680.668071441, 101779.825716651, 101998.733355457, 
    101779.585041833, 101384.053591, 101148.339135459, 101096.739349883, 
    101017.126636415, 100987.238807655, 100920.580424318, 100880.010074674, 
    100888.26119153, 101004.819082622, 101042.639363268, 101125.782349353, 
    101271.767323067, 101414.874544034, 101606.714170176, 101781.90582545, 
    101967.982450008, 102079.366590713, 102036.282211265, 101829.296739921,
  101498.647043559, 101590.9176954, 101617.915033384, 101637.802643964, 
    101648.185762942, 101655.587465239, 101658.006887633, 101549.42825388, 
    101414.618079725, 101373.424560394, 101351.03384233, 101279.222124666, 
    101130.397265545, 101055.783573411, 100985.0857455, 100980.935004011, 
    100935.286534163, 100896.981581297, 100779.214201905, 100638.338446691, 
    100455.513812383, 100365.634006852, 100280.18805953, 100314.217914751, 
    100429.553904417, 100663.751214393, 100811.813174929, 100901.524902021, 
    101010.647515613, 101164.233242571, 101286.631571935, 101379.069333755, 
    101445.325107445, 101498.821421146, 101521.036907936, 101495.177333539, 
    101475.52262969, 101380.590954348, 101245.617401119, 101122.593133959, 
    101083.032382908, 101027.109920763, 100965.681089336, 100868.736274192, 
    100845.638733495, 100806.63870496, 100789.709636642, 100730.892231111, 
    100731.226876586, 100656.195362061, 100620.062463698, 100541.660250164, 
    100462.584089641, 100519.284702863, 100618.483169607, 100730.59486643, 
    100851.037099314, 100994.659154739, 101129.958372846, 101331.846054031,
  101475.49557051, 101570.920009059, 101674.630218099, 101728.771159046, 
    101769.510444793, 101775.068660928, 101704.67979635, 101640.720658865, 
    101574.382411521, 101503.398083084, 101496.227909434, 101483.885943964, 
    101500.719290317, 101478.508725144, 101490.730004083, 101464.972200966, 
    101493.079514999, 101506.442828051, 101534.382393965, 101514.711231632, 
    101522.240678456, 101474.806810392, 101487.745795629, 101447.297047833, 
    101448.741711988, 101449.346100917, 101491.142897043, 101525.258984486, 
    101568.295073022, 101546.720496798, 101500.38695074, 101482.412130758, 
    101497.942828869, 101531.720763558, 101560.615239549, 101594.165172661, 
    101568.818695878, 101562.810678583, 101534.927138634, 101485.271491949, 
    101422.675613505, 101441.037784656, 101438.474919451, 101435.089671792, 
    101392.827173765, 101421.881442681, 101441.896959987, 101506.296721786, 
    101504.023500445, 101561.478585626, 101519.337418794, 101500.880468648, 
    101550.683255314, 101515.689136433, 101484.579866181, 101486.847559185, 
    101498.039007899, 101470.609948212, 101451.431054765, 101423.141133153 ;

 t =
  199.592302597963, 199.631103000267, 199.731954187836, 199.892616003787, 
    200.097555270638, 200.32094214551, 200.516784754057, 200.630608485976, 
    200.651370880938, 200.609578569847, 200.541354699461, 200.4600639894, 
    200.367096011648, 200.258081356635, 200.131678494282, 200.003927573354, 
    199.892093045302, 199.78951395173, 199.67327063218, 199.562612042923, 
    199.479736833425, 199.436427112334, 199.446431492281, 199.495730546513, 
    199.549832254666, 199.604520501067, 199.697689137597, 199.864710041022, 
    200.093779681868, 200.340566539804, 200.552259625836, 200.701276302059, 
    200.782756153405, 200.7833906832, 200.686856127812, 200.491170464732, 
    200.222261082732, 199.935938107253, 199.680606174414, 199.471038784987, 
    199.299652459908, 199.17323872267, 199.128354161206, 199.202004245832, 
    199.359077079051, 199.506090503528, 199.612484430338, 199.711922901369, 
    199.816793014736, 199.916139249983, 199.997437583028, 200.04825723153, 
    200.06355478738, 200.032336458477, 199.96631189711, 199.887308498887, 
    199.810491632393, 199.730691469998, 199.655116951929, 199.604483206791,
  199.925450534086, 199.981216668507, 200.13372177414, 200.374983049979, 
    200.666746595261, 200.968689298795, 201.213497199314, 201.320081014682, 
    201.28285515959, 201.159427975395, 201.016640981215, 200.883658495912, 
    200.771379174995, 200.674203060131, 200.572788065495, 200.477172369812, 
    200.407545496821, 200.338859718061, 200.224248971463, 200.078773906287, 
    199.945758232313, 199.862629278066, 199.864007266231, 199.931896031448, 
    200.010381034324, 200.095604476198, 200.236502900669, 200.462822228967, 
    200.753296999852, 201.044097788301, 201.25745758838, 201.374991871653, 
    201.427242945419, 201.406575723115, 201.277595633766, 201.023620969068, 
    200.67474741735, 200.313928085033, 200.00562786958, 199.761123711398, 
    199.573928575976, 199.465163976854, 199.478724977567, 199.645844456424, 
    199.924582984045, 200.192359977098, 200.373679113298, 200.483516015946, 
    200.545327071018, 200.577126788341, 200.591566679776, 200.576595520702, 
    200.535205988156, 200.455414739312, 200.357229008022, 200.262675215774, 
    200.183848343407, 200.096660938015, 200.004418550248, 199.940673718636,
  199.744781513231, 199.914256718427, 200.214409920574, 200.617360179337, 
    201.024747223831, 201.346435179694, 201.485950279302, 201.372767584886, 
    201.066836108378, 200.683142568019, 200.327292868912, 200.043685756443, 
    199.877844232157, 199.85781502703, 199.917492370117, 199.9983289047, 
    200.058369493754, 200.02806545364, 199.869574128922, 199.638192515119, 
    199.387877277734, 199.208849364091, 199.203422279425, 199.363656462519, 
    199.572566915159, 199.785805305591, 200.070728844411, 200.443013143122, 
    200.822614297206, 201.143713031253, 201.341847192701, 201.38421638141, 
    201.345298401764, 201.282948578685, 201.14389944696, 200.84584052779, 
    200.421451502179, 200.00681344595, 199.656631388896, 199.360541466825, 
    199.14599754243, 199.085672435604, 199.226941252801, 199.564065741742, 
    200.023699867917, 200.448535551099, 200.717131468681, 200.801164827762, 
    200.709143038557, 200.510624205462, 200.310857959432, 200.123534038996, 
    199.985918823302, 199.870278463294, 199.810564689902, 199.802795120091, 
    199.809558043709, 199.777525661617, 199.711729725736, 199.683753027175,
  198.813626070185, 199.158986036996, 199.627864744577, 200.160256266574, 
    200.623623253207, 200.864117088923, 200.781735620651, 200.390995226515, 
    199.824482274509, 199.223765018052, 198.69225842097, 198.246625464903, 
    197.991561721856, 198.105138108831, 198.488106862037, 198.875209917554, 
    199.041959326812, 198.902255067274, 198.524256150457, 198.120422776864, 
    197.754283879839, 197.52804051378, 197.557076137182, 197.838677763684, 
    198.228311776218, 198.64866693467, 199.141249850207, 199.671836733273, 
    200.066037593716, 200.26086896737, 200.335026610284, 200.27629681715, 
    200.145458434459, 200.058740328064, 199.982932145149, 199.734988702051, 
    199.342332480579, 198.978689763372, 198.64265554624, 198.322820390541, 
    198.141459621883, 198.230337302711, 198.595370204332, 199.122716273707, 
    199.641829159866, 199.98647687541, 200.106596249157, 200.023669500759, 
    199.71862786998, 199.269902761839, 198.872993350988, 198.549303124569, 
    198.402247374352, 198.389745298667, 198.520267551177, 198.727735192993, 
    198.820080794775, 198.772285728007, 198.671469694149, 198.647026352616,
  198.27177169786, 198.742255912744, 199.315734313932, 199.897371339361, 
    200.359948915917, 200.535691314823, 200.35927551603, 199.924949090263, 
    199.330086169064, 198.665856285035, 198.042667303558, 197.482635890829, 
    197.119520606414, 197.266701392985, 197.835195092286, 198.339553763094, 
    198.478815953183, 198.22439010637, 197.650427994835, 197.067516663093, 
    196.641410409783, 196.481794550396, 196.629327985159, 197.039139885895, 
    197.582657417974, 198.18477677987, 198.804275829209, 199.362413123988, 
    199.653029088601, 199.576374980457, 199.317720083802, 199.03686382968, 
    198.89995519903, 198.950655967047, 199.063529863595, 198.990505226734, 
    198.75355662612, 198.500929788027, 198.208223031476, 197.938423894621, 
    197.885803160602, 198.139155318154, 198.615513384798, 199.131104917232, 
    199.510955642597, 199.659024904865, 199.580116095284, 199.333081499491, 
    198.916549920377, 198.433254494224, 198.05605526358, 197.713977419289, 
    197.562858694346, 197.648783925538, 197.92635060358, 198.262190792517, 
    198.337240530356, 198.203194194284, 198.058390816553, 198.034817661849,
  198.937766800522, 199.378862901994, 199.924167284663, 200.441900343408, 
    200.827224031058, 200.990625476238, 200.897309110033, 200.618864003997, 
    200.181564650821, 199.613998887189, 198.983091583902, 198.347030011959, 
    197.856354212493, 197.870456627708, 198.431509424617, 198.97692508607, 
    199.135205071391, 198.873711540888, 198.238990745813, 197.579817494844, 
    197.172597878355, 197.088718428204, 197.353762305792, 197.89826630309, 
    198.564087596207, 199.248896670098, 199.861576972738, 200.25445850994, 
    200.212422489697, 199.775398283844, 199.153661619413, 198.657419145184, 
    198.616608196145, 198.978344443701, 199.371695654673, 199.518116209905, 
    199.425895663568, 199.218774286518, 198.944338234565, 198.750162861572, 
    198.807293796669, 199.126797161784, 199.590707523985, 200.01113682887, 
    200.236675555464, 200.213934135267, 199.968933435599, 199.597738976311, 
    199.166919297141, 198.80613007738, 198.561749801842, 198.310183827336, 
    198.209165549116, 198.396376260841, 198.756180625289, 199.008102754839, 
    198.971509894537, 198.817890375389, 198.71624809131, 198.718856697764,
  199.468938785267, 199.746343042481, 200.264885640233, 200.799307962387, 
    201.187287972447, 201.364687823852, 201.345163759808, 201.220378142663, 
    200.97932418323, 200.594250421451, 200.052751072066, 199.422214940597, 
    198.841924275609, 198.642398630235, 199.050269137882, 199.669323207652, 
    200.028156686643, 199.896274809802, 199.320690987659, 198.647441033344, 
    198.165872236427, 197.964443275584, 198.191936305371, 198.832089684652, 
    199.66059838197, 200.451219513806, 201.004151536921, 201.167557397172, 
    200.814529868517, 200.148624018046, 199.383120991314, 198.942875215344, 
    199.10824731445, 199.672579767983, 200.084759895193, 200.167771094173, 
    200.048559955598, 199.894763241948, 199.724712360714, 199.612023496662, 
    199.667017008079, 199.927888948017, 200.330942504098, 200.713413442935, 
    200.903819251949, 200.783835877041, 200.374816063361, 199.841531051172, 
    199.370642946036, 199.155395223596, 199.122641487494, 199.065805967836, 
    199.004343588847, 199.137833233884, 199.538339084755, 199.870585152783, 
    199.958157705803, 199.880438792344, 199.701546365556, 199.494348467994,
  198.448112855695, 198.354611013293, 198.728868336993, 199.316380836934, 
    199.79403116714, 200.005499925149, 199.986681621127, 199.959375733492, 
    199.916472122982, 199.742737462745, 199.386100288375, 198.895591537667, 
    198.365829775093, 198.004132576714, 198.061450403236, 198.512771018877, 
    199.123932187329, 199.430874598043, 199.211486449103, 198.613405452253, 
    197.929414433977, 197.40356151974, 197.327965358493, 197.871397861698, 
    198.835639679273, 199.725297830638, 200.085368082906, 199.928953443704, 
    199.386031776095, 198.761776597613, 198.266743904794, 198.170096710373, 
    198.41391650884, 198.774680929286, 198.886267152027, 198.743207447002, 
    198.609154244075, 198.681026842838, 198.846271254613, 198.944125173226, 
    198.942818972897, 198.966709387328, 199.149155931741, 199.505726712438, 
    199.844168672597, 199.85140388845, 199.45483469524, 198.809580467374, 
    198.167797788754, 197.859611842392, 197.936977186745, 198.163259504691, 
    198.218548157533, 198.115014051873, 198.1926679382, 198.557752668518, 
    199.061087852164, 199.366370956955, 199.261747362555, 198.84460292621,
  197.485930857678, 197.019818372692, 197.201895561925, 197.805867406745, 
    198.350370518934, 198.583615055967, 198.478395457053, 198.407310549954, 
    198.450691963437, 198.439158293822, 198.294734348496, 197.997424250824, 
    197.615467503654, 197.255442031252, 197.102529470095, 197.311811051274, 
    197.910422679403, 198.566184591881, 198.81770599644, 198.468817940017, 
    197.724338140697, 196.932991398967, 196.470632589878, 196.715726910412, 
    197.667118273752, 198.570347547162, 198.71122967919, 198.221418635834, 
    197.430221844445, 196.808140980382, 196.687634903507, 197.099568018172, 
    197.579347149138, 197.825720124614, 197.684919362109, 197.28817327461, 
    196.99979888361, 197.130125348385, 197.614586291391, 198.054621237893, 
    198.133785793687, 197.953725042329, 197.830236454786, 198.056196080487, 
    198.536103308907, 198.780904128645, 198.57011209624, 197.965907355598, 
    197.227821256842, 196.76451533989, 196.770352581149, 197.088045611668, 
    197.205666419854, 196.943229549179, 196.598121652703, 196.623097357434, 
    197.265132242531, 198.08254785051, 198.422861021731, 198.114028385677,
  197.5134829456, 196.944617330308, 197.046071825314, 197.62502348085, 
    198.161844347888, 198.368966236773, 198.173531381369, 198.018783271948, 
    198.061430667878, 198.131590257702, 198.122379709768, 197.921446982702, 
    197.619936793757, 197.323568470083, 197.152715436221, 197.285048638712, 
    197.822753961333, 198.569172895512, 199.007248056168, 198.844079816698, 
    198.16595031969, 197.314536253415, 196.730018868748, 196.844187956897, 
    197.72913335811, 198.475588226684, 198.454427766617, 197.801336310951, 
    196.85090861976, 196.20593400157, 196.280422982296, 196.977580932572, 
    197.680530000096, 197.997569172916, 197.806564556565, 197.31204925314, 
    196.902648128082, 196.994797825051, 197.584353315729, 198.160576501024, 
    198.284328642877, 198.010801157452, 197.694140964105, 197.764900474119, 
    198.25282328335, 198.655964724116, 198.65227811331, 198.181742441883, 
    197.476943605846, 196.968619353371, 196.935358254191, 197.224878909066, 
    197.288545612313, 196.956882630364, 196.394991024497, 196.117522272038, 
    196.658334362852, 197.680111197301, 198.298723643018, 198.154816315995,
  198.166109085876, 197.718670143435, 197.86168227072, 198.369607608057, 
    198.793450206587, 198.908504936618, 198.690993492582, 198.512396667806, 
    198.566541502908, 198.67011073685, 198.66255442265, 198.424151351069, 
    198.117772276422, 197.891735389794, 197.849998798018, 198.10665993907, 
    198.677352006052, 199.297136934201, 199.565704814004, 199.314718369792, 
    198.690725808071, 198.035269907306, 197.68129614681, 197.93520103824, 
    198.722931139366, 199.179410889798, 199.042652872112, 198.371641439503, 
    197.476189927944, 196.950977014733, 197.080876424779, 197.7319570849, 
    198.397313053343, 198.7212284182, 198.5805281666, 198.208118865396, 
    197.863282454832, 197.963307975476, 198.511882923795, 199.005063445837, 
    199.075262984366, 198.754841079178, 198.390987981186, 198.401463363339, 
    198.77139605576, 199.120481880218, 199.158232177865, 198.818050246871, 
    198.316276705667, 197.956185781121, 197.987116929256, 198.223657072334, 
    198.187964808669, 197.833057589277, 197.246013805985, 196.931446448565, 
    197.40217386718, 198.309189620928, 198.838359180219, 198.723822600565,
  199.641955409729, 199.431669295405, 199.670215080691, 200.063453434526, 
    200.291822159985, 200.229512907391, 200.018076015997, 199.891370308544, 
    199.98823486655, 200.056917508163, 199.974392905842, 199.676282742029, 
    199.396510789061, 199.324214877096, 199.545065181078, 200.032738777083, 
    200.587110551674, 200.84423935639, 200.780242526822, 200.386860036893, 
    199.868432218779, 199.591695869976, 199.618184911359, 200.035059503488, 
    200.578885970644, 200.670005940932, 200.424434628647, 199.853721051106, 
    199.202883004278, 198.956638029292, 199.156376634439, 199.579947395386, 
    199.972684533674, 200.183496369922, 200.077062289701, 199.875609449205, 
    199.718992210914, 199.890333068829, 200.336224521985, 200.636983405007, 
    200.605632519331, 200.296665053459, 199.991350344062, 199.992817812916, 
    200.163951929184, 200.2945713224, 200.240193398709, 200.001834516286, 
    199.762256009081, 199.65534366822, 199.78956330339, 199.952345481649, 
    199.825002417001, 199.49596919313, 199.043589284655, 198.920122405191, 
    199.394323032761, 200.010122477167, 200.234707331376, 200.056809522668,
  200.473296344829, 200.441424752327, 200.678958349945, 200.918516462326, 
    200.956552022289, 200.723091611172, 200.525940020957, 200.472508457677, 
    200.597371060414, 200.593157561086, 200.474003063485, 200.253130275181, 
    200.147547411406, 200.296157360971, 200.693653157222, 201.208414708891, 
    201.559490813672, 201.537219487268, 201.316024304306, 200.882014152838, 
    200.457138758545, 200.50571123716, 200.831560678168, 201.22579454473, 
    201.397276457415, 201.232054205466, 201.003522505839, 200.657457121342, 
    200.253185454957, 200.154639454359, 200.362553394409, 200.604148733558, 
    200.765528887011, 200.872139048546, 200.802617853893, 200.723083041081, 
    200.731974781426, 200.902646174949, 201.160028006192, 201.277512234295, 
    201.204036684047, 200.970540553361, 200.735983962232, 200.703512138846, 
    200.748936469414, 200.752492313878, 200.670067358296, 200.520078028079, 
    200.450192550345, 200.519108630864, 200.672244639888, 200.731752862692, 
    200.587200372453, 200.364686349462, 200.104714472775, 200.10985779648, 
    200.465145414594, 200.803151432196, 200.827806544744, 200.682191054799,
  201.213225510545, 201.166835543629, 201.270714839611, 201.37550537134, 
    201.324990086747, 201.082379320499, 200.962481306926, 200.995956365887, 
    201.095973310753, 201.017526279202, 200.891099818738, 200.813033119912, 
    200.865724272731, 201.079500872488, 201.395316575206, 201.681516167276, 
    201.76670295158, 201.757393321422, 201.692231811594, 201.40827235103, 
    201.075956075215, 201.189995122758, 201.557166511341, 201.81492663249, 
    201.746759931066, 201.570017408439, 201.47269399979, 201.328677087196, 
    201.125151299054, 201.055029029273, 201.188090739647, 201.31703109918, 
    201.35013936096, 201.369651479787, 201.321315159999, 201.287934158944, 
    201.349721325709, 201.47663855592, 201.609607336194, 201.647923717432, 
    201.571079750039, 201.36274141706, 201.168463850806, 201.156910392398, 
    201.202814218407, 201.20117036627, 201.18331549404, 201.127720965669, 
    201.108346069018, 201.173613329739, 201.223083981493, 201.16065459979, 
    201.079743557461, 201.038714778534, 200.94457273968, 200.937378451857, 
    201.093228584694, 201.285737192623, 201.319924072079, 201.296636239629,
  202.281128399983, 202.174317384615, 202.183902282345, 202.196135777651, 
    202.089228467659, 201.946467982868, 201.939131149378, 202.047091741652, 
    202.150160623985, 202.131660791028, 202.004701967929, 201.929182231624, 
    201.93459873504, 202.027913871461, 202.17850666923, 202.292775710951, 
    202.295938725162, 202.40040339815, 202.492591335442, 202.422978333309, 
    202.266666952811, 202.298371892207, 202.475203686205, 202.593449698724, 
    202.486915616929, 202.407280373555, 202.418866882487, 202.398256235396, 
    202.399756349372, 202.37264124627, 202.399210244757, 202.401295541644, 
    202.3114410158, 202.232821203222, 202.191752199712, 202.19277899535, 
    202.267398417301, 202.391431505571, 202.515532414131, 202.539412611326, 
    202.465954562056, 202.318811656422, 202.240022548479, 202.297290346244, 
    202.317551796671, 202.256173931376, 202.220798534059, 202.171503678984, 
    202.150285293746, 202.201814576557, 202.183544018307, 202.011884222124, 
    201.959863852426, 202.041740696822, 202.056502837546, 202.032604839674, 
    202.07407065357, 202.222871000044, 202.358430896211, 202.414399487383,
  202.386516519161, 202.267030767596, 202.378273066683, 202.433008545321, 
    202.347394948355, 202.349805373492, 202.448279893784, 202.631049610784, 
    202.827361753103, 202.874316929906, 202.669053832267, 202.492135754915, 
    202.409415422156, 202.422620106113, 202.501927380974, 202.552975255795, 
    202.533541984178, 202.569576423265, 202.56117823678, 202.539935320285, 
    202.520947357138, 202.552469465724, 202.620265993283, 202.674370717175, 
    202.569923878364, 202.510390647561, 202.541104878651, 202.581706643803, 
    202.689332310414, 202.6892441831, 202.66916514168, 202.614276720316, 
    202.47365472681, 202.336160185186, 202.28527670572, 202.311285294881, 
    202.392266489274, 202.542076139595, 202.726730639659, 202.790019717988, 
    202.722561395316, 202.609789063794, 202.55770098193, 202.562571664569, 
    202.497193469629, 202.415414918844, 202.406393221663, 202.378392740735, 
    202.369165519715, 202.420992607534, 202.392358940459, 202.196524439297, 
    202.130920806496, 202.207092624452, 202.265923810763, 202.273893555593, 
    202.291904065293, 202.425980200592, 202.689171477895, 202.763829093729,
  201.105874470791, 201.100406974456, 201.304475401087, 201.312268793347, 
    201.143074728591, 201.098131592507, 201.120851793788, 201.267279389605, 
    201.562668172102, 201.779931434368, 201.780627457301, 201.69059514426, 
    201.577244544257, 201.516684463659, 201.508651367797, 201.485053452921, 
    201.46118383068, 201.466399046118, 201.407989930795, 201.382955438949, 
    201.38521694024, 201.454277056699, 201.540505008593, 201.555927231927, 
    201.375433672908, 201.218119197833, 201.19784543263, 201.295666775342, 
    201.490543698467, 201.59693764053, 201.647057234143, 201.579829538758, 
    201.428484001518, 201.240934751399, 201.127926290216, 201.132320301533, 
    201.193096487911, 201.344183945922, 201.56545304613, 201.674803851175, 
    201.6316049083, 201.500875996819, 201.370252773686, 201.286143050101, 
    201.238226725847, 201.298383416386, 201.408901089709, 201.412828942136, 
    201.352636482984, 201.274948494925, 201.176520349776, 201.048394695858, 
    201.020782354372, 201.040590737723, 201.050091755113, 201.049191850238, 
    201.073625314884, 201.169042997751, 201.451596197436, 201.544358138887,
  200.457208020337, 200.600627775773, 200.766445085137, 200.658695042864, 
    200.379501992268, 200.193506888721, 200.159959051097, 200.417920530747, 
    200.881492064797, 201.158314717164, 201.185079926141, 201.052599033083, 
    200.912278077891, 200.826400220702, 200.745363986095, 200.644201348986, 
    200.621331534948, 200.670081702674, 200.634010510041, 200.57519712089, 
    200.537473759589, 200.668670498033, 200.855042651151, 200.850338930202, 
    200.564184196878, 200.26841305199, 200.153083417943, 200.265131602254, 
    200.562861149189, 200.91898622909, 201.262053214654, 201.293252570222, 
    201.048704338528, 200.619896243786, 200.289829022617, 200.230648433139, 
    200.336307776342, 200.615867228439, 200.978592412832, 201.151128388213, 
    201.06018709287, 200.772139831747, 200.439274423229, 200.215103174651, 
    200.214000730343, 200.477371906456, 200.762592440744, 200.820520583299, 
    200.718859121984, 200.529592256917, 200.334051442783, 200.1976241956, 
    200.1567040591, 200.14207121777, 200.132612485116, 200.195054606259, 
    200.344963296675, 200.442882819041, 200.626470402943, 200.688840294464,
  200.025483430949, 200.16208883287, 200.313588748616, 200.213688182892, 
    199.913595102692, 199.578945078437, 199.457159567169, 199.837498014033, 
    200.589263318679, 201.039711065693, 201.012585788289, 200.648141762678, 
    200.273131591484, 200.097802170007, 200.054831651363, 200.044432329585, 
    200.102085232929, 200.195405788936, 200.160924644118, 200.038915629557, 
    199.916144055078, 200.079124573273, 200.367134834657, 200.411516440404, 
    200.134086471815, 199.790609936755, 199.62840687339, 199.728355779226, 
    200.048032676646, 200.504469872656, 201.036196596741, 201.238698672334, 
    200.985033674728, 200.320989492277, 199.680506629958, 199.407286593517, 
    199.463090763364, 199.919203575643, 200.599348362119, 201.013906220406, 
    200.959187102964, 200.499767817349, 199.883859695177, 199.41997174576, 
    199.340501041543, 199.679936618532, 200.144417395864, 200.372293549977, 
    200.376297420661, 200.221448294299, 199.975937237797, 199.739637238205, 
    199.573253617133, 199.482002551712, 199.458807211945, 199.662248641179, 
    200.080451213873, 200.317721543376, 200.394403633302, 200.243350533172,
  198.793407369955, 198.789017315693, 198.904292936824, 198.815824252696, 
    198.495882684834, 198.008478868489, 197.715295378614, 198.048286658139, 
    199.034194857732, 199.804116024622, 199.863316118556, 199.322511698704, 
    198.564555658753, 198.130267186998, 198.214466779197, 198.620047714388, 
    199.003291040746, 199.12920558678, 198.939536007096, 198.634278790921, 
    198.422185184682, 198.646306495756, 199.004286128174, 199.099073335961, 
    198.889156737865, 198.546163685228, 198.365896567428, 198.448978172239, 
    198.756197741766, 199.223797691081, 199.827895879143, 200.210498988022, 
    200.027828598842, 199.255370438114, 198.305435802773, 197.601225043893, 
    197.345365719658, 197.840319194022, 198.882186376654, 199.694423752905, 
    199.826621632831, 199.31781668854, 198.474553418244, 197.742364960171, 
    197.469627758775, 197.758017180375, 198.409942614757, 198.98336969176, 
    199.298780373215, 199.302239468507, 199.040595330121, 198.653688069122, 
    198.243554048026, 197.9377903084, 197.80783043139, 198.063400210034, 
    198.693135810417, 199.184504322592, 199.335127001616, 199.113968919495,
  198.221704432865, 198.148506305094, 198.205050154027, 198.013097013938, 
    197.539633153928, 196.849673610595, 196.334807195508, 196.533836294342, 
    197.642709038047, 198.693594051791, 198.854871373202, 198.211458363155, 
    197.162500404924, 196.468372290433, 196.675366563475, 197.582272798516, 
    198.400163183235, 198.611071666639, 198.241204377327, 197.695950454543, 
    197.377636018492, 197.6448646534, 198.085850918047, 198.235251613086, 
    198.034649097847, 197.588365548619, 197.279834838421, 197.351544608965, 
    197.753649740072, 198.335099296068, 199.036322336768, 199.564463145478, 
    199.432841323671, 198.598687407314, 197.453743242996, 196.421391648673, 
    195.903353846926, 196.396124609721, 197.648174115494, 198.708648439145, 
    198.947977723217, 198.400474668592, 197.422099467524, 196.521148254654, 
    196.103106473721, 196.368001370275, 197.203807165087, 198.102800907396, 
    198.699799081932, 198.867802373005, 198.661471438684, 198.205189016116, 
    197.616845313813, 197.07106617434, 196.701708097593, 196.794169022806, 
    197.430803098791, 198.160314033553, 198.528415308627, 198.490707039997,
  198.905702879998, 198.738136377768, 198.613804463776, 198.226709598317, 
    197.597394605101, 196.861360985921, 196.342172243993, 196.543197341785, 
    197.604251929708, 198.566522282061, 198.612577634039, 197.883144750032, 
    196.821343717449, 196.183431256679, 196.577755929701, 197.748455047779, 
    198.751654537677, 199.003051214735, 198.591100771163, 197.991726261388, 
    197.650258353922, 197.871702346101, 198.263977124647, 198.312614950729, 
    198.018442923194, 197.488490192782, 197.091610662671, 197.206971302572, 
    197.764783042513, 198.508059655596, 199.2772086787, 199.763075521379, 
    199.54296860815, 198.67045658231, 197.554135264445, 196.567888928647, 
    196.160391392102, 196.763249480626, 197.949691304552, 198.845735933519, 
    198.928508306334, 198.300914607485, 197.323611181691, 196.45854393356, 
    196.102870918749, 196.509901689766, 197.480545100735, 198.442070117891, 
    199.065283184618, 199.259051952296, 199.088315896478, 198.626312565053, 
    197.963036596952, 197.25333848771, 196.647276031209, 196.54265825896, 
    197.157970301143, 198.135536397283, 198.837259866507, 199.078046102662,
  199.748686826344, 199.27778362655, 198.895353036917, 198.468684976879, 
    197.950914905868, 197.470716295197, 197.256535798763, 197.587299145965, 
    198.413626251024, 198.963879920237, 198.744498143694, 198.022499808208, 
    197.265828623102, 197.025754304726, 197.644096805373, 198.763418388169, 
    199.616119773958, 199.791137713501, 199.416787390728, 198.901569342749, 
    198.546835407943, 198.526698700786, 198.60752753218, 198.418287351064, 
    198.060977343818, 197.620683187014, 197.35909651458, 197.618614399286, 
    198.289062384969, 199.078551099742, 199.743381893889, 200.01438191863, 
    199.698603256515, 198.946744193281, 198.127702903355, 197.568238693356, 
    197.598045009421, 198.279360568835, 199.05915077239, 199.427625208044, 
    199.181371546663, 198.470198316339, 197.617314753671, 196.991152962905, 
    196.900914299691, 197.490642065525, 198.396135446458, 199.071604497419, 
    199.444106613956, 199.557939824348, 199.39190234454, 198.942192820278, 
    198.307578484637, 197.623785024728, 196.995571588184, 196.829800056189, 
    197.449032433194, 198.59669332296, 199.581667984863, 199.994678428791,
  200.187773471693, 199.557720394685, 199.235729652164, 199.070652084612, 
    198.854039702492, 198.769404371782, 198.979443417092, 199.3266764035, 
    199.64286620581, 199.674688259513, 199.314692534306, 198.821908340682, 
    198.541295809677, 198.735770563891, 199.423172574944, 200.253650111218, 
    200.778222412623, 200.799441991581, 200.444304814849, 199.981775630426, 
    199.523214012252, 199.133053396801, 198.852995270112, 198.583728548467, 
    198.386698785655, 198.262261584952, 198.311393023357, 198.682662636759, 
    199.277569921611, 199.886606569575, 200.319984116121, 200.42955050266, 
    200.182252880161, 199.786978398504, 199.53194688739, 199.567389851748, 
    199.892015112085, 200.273918676104, 200.419038592148, 200.198841496834, 
    199.646265661263, 198.888900496761, 198.235484423046, 197.984496635759, 
    198.229234260917, 198.82013922824, 199.331455388365, 199.455093241226, 
    199.488592468736, 199.68690678624, 199.724655145764, 199.40506796936, 
    198.876470297172, 198.303317398924, 197.817844339452, 197.74178639462, 
    198.291461196874, 199.296576709642, 200.208368919365, 200.552300800139,
  200.088893253039, 199.548292267843, 199.356641782753, 199.402446204426, 
    199.470527191872, 199.65298386703, 199.977318009437, 200.170458705907, 
    200.138889178331, 199.941004138127, 199.623645714064, 199.400249828807, 
    199.440334932923, 199.796997237617, 200.355721453897, 200.838039244748, 
    201.030259713147, 200.871971259787, 200.458090357353, 199.935184834046, 
    199.366326152042, 198.835369275314, 198.525846247017, 198.461707883348, 
    198.547543996739, 198.709571593396, 198.98956432621, 199.403416757117, 
    199.851753400366, 200.215210527421, 200.419573373203, 200.438987900915, 
    200.343685887155, 200.322658635607, 200.49680159455, 200.81524409789, 
    201.06616648875, 201.012269368143, 200.714356047539, 200.155458175476, 
    199.46064866819, 198.8125502932, 198.500814466291, 198.59490291881, 
    198.898088049482, 199.186662677498, 199.264894911019, 199.072273851087, 
    198.990545700138, 199.358253558878, 199.666118568762, 199.587301995179, 
    199.280270729975, 198.932512050275, 198.65404251086, 198.620336243918, 
    198.935929165386, 199.551770943114, 200.156627443202, 200.405844334092,
  199.672687015645, 199.339465822255, 199.174377451439, 199.208979460959, 
    199.382291687595, 199.685923357783, 199.991210902835, 200.099800254538, 
    200.005065026363, 199.794268081768, 199.526034053772, 199.389450686464, 
    199.477207094757, 199.769609806221, 200.144237090792, 200.381831349755, 
    200.372238222555, 200.102451305332, 199.644633254532, 199.108673684973, 
    198.556259861019, 198.11725745431, 197.92256156203, 197.982163336143, 
    198.213826014132, 198.549350231965, 198.958893887917, 199.385421798674, 
    199.755817435057, 200.0165120883, 200.14527899575, 200.182785764376, 
    200.208645802587, 200.278005378702, 200.458601503633, 200.747245075818, 
    200.877140695159, 200.592634977004, 200.084270168955, 199.380009378005, 
    198.651450545581, 198.151387053296, 198.045866371994, 198.202887764545, 
    198.417868308159, 198.581172029478, 198.633325488976, 198.552252187611, 
    198.488480439262, 198.692849285014, 198.972857703249, 199.113422906924, 
    199.104413126486, 198.989393755147, 198.863445331237, 198.871619392842, 
    199.05601502309, 199.372804189126, 199.667214807037, 199.837999534726,
  199.528577019934, 199.372328554741, 199.219255608941, 199.181174953061, 
    199.317772524265, 199.594571234405, 199.838696964916, 199.932207161942, 
    199.905701026384, 199.807690567105, 199.634257382221, 199.478539330645, 
    199.445720085212, 199.574856739142, 199.781791750333, 199.895475994151, 
    199.828921664597, 199.560103893746, 199.108712898402, 198.602286364023, 
    198.136174000588, 197.810600389175, 197.65646262947, 197.675058604625, 
    197.871768137081, 198.220658718832, 198.652234853298, 199.084188327866, 
    199.467633249614, 199.766624716516, 199.954339826767, 200.059567083605, 
    200.133779341625, 200.191034943094, 200.296674583153, 200.47543202185, 
    200.532203533176, 200.256344227993, 199.747674414816, 199.072770558125, 
    198.383004828485, 197.886509098768, 197.666326148207, 197.665249670721, 
    197.813481807783, 198.002685781874, 198.151820080209, 198.227674286913, 
    198.248837381842, 198.339114953752, 198.498871312887, 198.628206411758, 
    198.72272650249, 198.774672679998, 198.832670572642, 198.957968430551, 
    199.123423919216, 199.300243175253, 199.43879711417, 199.559413990189,
  199.563276840686, 199.5522915196, 199.47998544867, 199.417818470489, 
    199.446999729066, 199.581507224339, 199.737654813664, 199.833163318563, 
    199.845075194212, 199.795466188751, 199.700627898087, 199.59683259565, 
    199.525796962369, 199.50082970616, 199.488693505057, 199.445943085924, 
    199.349730635173, 199.17519308442, 198.876787942237, 198.513574919775, 
    198.149387221562, 197.840999813482, 197.627271367646, 197.559549529766, 
    197.668022765168, 197.925767343833, 198.267312100976, 198.640681702791, 
    199.024447350664, 199.370552776363, 199.617054991639, 199.766535336821, 
    199.871913674194, 199.969021841662, 200.085497705293, 200.213292782578, 
    200.278434443729, 200.184408630195, 199.908468458637, 199.4716320612, 
    198.964026024853, 198.540832766649, 198.263663299724, 198.123718276166, 
    198.067153592188, 198.017208056177, 197.980992450428, 197.98132422998, 
    198.011515397882, 198.079600686078, 198.14907558945, 198.191094916103, 
    198.2753526549, 198.422322297996, 198.621465940566, 198.838495055261, 
    199.038415085385, 199.217908373215, 199.361116652052, 199.490733842502,
  199.775980560716, 199.826624087702, 199.841035966137, 199.848740895578, 
    199.883214543563, 199.952415883452, 200.025036671968, 200.062157495331, 
    200.047954450696, 199.997297210152, 199.925240070427, 199.837823762514, 
    199.740778520753, 199.641158943761, 199.546007596529, 199.472066942666, 
    199.41121013987, 199.335200566612, 199.193460572359, 198.990450982689, 
    198.750882001109, 198.51109152544, 198.314639876566, 198.214985959892, 
    198.235447302199, 198.354596983364, 198.534190198528, 198.747035502699, 
    198.972887080861, 199.173781776681, 199.331694422277, 199.483053685455, 
    199.669481456939, 199.892844500556, 200.126831270649, 200.334453618466, 
    200.481599771775, 200.525235541313, 200.418154324323, 200.156350551711, 
    199.801364425044, 199.458602101623, 199.171055003088, 198.940400732437, 
    198.743249448746, 198.568817553593, 198.447470529527, 198.381793227975, 
    198.343109005189, 198.316167709471, 198.285223573377, 198.270811750809, 
    198.324486589019, 198.458581214609, 198.645553480285, 198.851328780692, 
    199.07694591123, 199.31289043773, 199.516363564806, 199.672765905304,
  199.505471640925, 199.573607216816, 199.628179558444, 199.679131836719, 
    199.73372238768, 199.791348393886, 199.835663376628, 199.850383518591, 
    199.834861016832, 199.79825953169, 199.745484073017, 199.676249995665, 
    199.595193987988, 199.51362655912, 199.444609026659, 199.404554714496, 
    199.38123925889, 199.352748417998, 199.286792110154, 199.173854598935, 
    199.023695635941, 198.86124427138, 198.715633252667, 198.620923669143, 
    198.594343737474, 198.624337853433, 198.689285509629, 198.769492182293, 
    198.845252160134, 198.899211928843, 198.95500540275, 199.067081895793, 
    199.262859125221, 199.523685504689, 199.805442725795, 200.060598579508, 
    200.251435133846, 200.340824165221, 200.291119459226, 200.100651686881, 
    199.825596737399, 199.539648563239, 199.276310663554, 199.043498856462, 
    198.84000982517, 198.674658311647, 198.559906851335, 198.483816741808, 
    198.421892961603, 198.366992865926, 198.326222545709, 198.320955878866, 
    198.370612772237, 198.475632949975, 198.612988709, 198.763519318843, 
    198.937246170728, 199.123194401409, 199.285685038358, 199.412233586054,
  212.299979432734, 212.06781029898, 211.855761765126, 211.748125242497, 
    211.763221995897, 212.12257479035, 212.527972829108, 212.441324714399, 
    212.218119073442, 212.085381261847, 212.044187386995, 212.002233488866, 
    212.026405101432, 212.122426770759, 212.315651949914, 212.560158246042, 
    212.759772546615, 212.83327989901, 212.635198579076, 212.579004298353, 
    212.752403220248, 212.948713945108, 212.720810843382, 212.10109282435, 
    211.830531141047, 211.967035312759, 212.355995900599, 212.514858832208, 
    211.846145645237, 211.207664895124, 210.95948666351, 210.777756058136, 
    210.819641832912, 211.140182823984, 211.552556319266, 211.924758084126, 
    212.284632745419, 212.577958759283, 212.843380360362, 213.102021384984, 
    213.388804423794, 213.553083209213, 213.640720982491, 213.747199130268, 
    213.685738015393, 213.318111386255, 212.887584960631, 212.582134537692, 
    212.459994820807, 212.383281490497, 212.300216765818, 212.306603130447, 
    212.402641479169, 212.500910425891, 212.699861547704, 212.742127600686, 
    212.6865352048, 212.676025957727, 212.711663871663, 212.513852102495,
  214.497151419508, 213.977357446485, 213.508783731028, 212.963821178042, 
    212.500457743552, 211.920620604982, 211.49309603927, 211.514504601478, 
    211.721232729647, 212.105552530266, 212.611535451222, 213.219897163857, 
    213.76768077524, 214.299261769899, 214.576925432378, 214.812782360487, 
    214.927351043233, 215.213582600175, 215.773772020066, 216.014741082582, 
    216.061606291433, 216.186692579083, 216.387298720466, 216.671783478429, 
    216.852584787981, 217.244875895593, 217.219117518403, 216.455214672446, 
    216.282977649656, 216.012244366936, 215.244185282641, 214.783458471721, 
    214.741336015231, 214.742940575343, 214.838359665979, 215.162102870675, 
    215.555975920051, 215.822522029634, 215.911323912162, 215.848900440489, 
    215.73356227059, 215.798987424043, 215.612947994145, 214.524087522498, 
    213.681808962539, 214.208731839748, 214.770768689681, 214.539889106084, 
    214.086318412745, 213.98818435472, 214.181097073179, 214.282901644277, 
    214.25061499428, 214.397566695256, 214.490524467729, 214.717088400921, 
    215.019238224473, 215.112906064012, 215.002473912384, 214.85425502345,
  213.582263826266, 212.256780413113, 211.078298467575, 210.727869840636, 
    210.65774032221, 210.95344737243, 211.504587816813, 212.568238996364, 
    214.101850561698, 215.193719296042, 215.444223367709, 215.406370756275, 
    215.461567276815, 215.593539679379, 216.158321670634, 216.553902302768, 
    216.967774472619, 216.920514141613, 217.419515690462, 217.336499335835, 
    216.982511205879, 216.856954083359, 216.473437063932, 216.15532762456, 
    216.804860156702, 217.16562778026, 217.82731505218, 218.847589707034, 
    218.0352766581, 217.255552228996, 217.668087631078, 217.620285337906, 
    217.175260776534, 217.554892822657, 218.374584340543, 219.10583976754, 
    219.839657295706, 220.356640037396, 220.101211592129, 218.979298623829, 
    217.560069105645, 215.949771177044, 214.64803238982, 213.993240895811, 
    212.96376750895, 212.0342396814, 212.856904565332, 214.637747563097, 
    216.328649689333, 217.32242201322, 217.617647033154, 217.719191345667, 
    217.615187237398, 217.523657615679, 217.950827211554, 218.053932047113, 
    217.386241667545, 216.708258746571, 215.992612006214, 214.886979892126,
  212.667168964723, 212.85393720424, 213.570452486422, 214.095039259794, 
    215.49518918329, 216.410391385443, 217.134948752383, 218.285676534147, 
    218.147571254928, 217.163145524981, 216.096888875451, 215.600843193118, 
    215.140045629146, 214.441033318532, 214.123497361284, 215.567395577976, 
    216.646601702513, 218.248121329369, 218.101381229466, 217.242264399979, 
    216.522803547047, 216.320488407572, 215.976684045793, 215.749380124998, 
    215.185739459463, 215.909866276403, 216.373364313196, 216.394736728967, 
    217.931514129965, 217.289994459314, 215.639510703103, 216.672342195904, 
    218.28957295573, 219.501915829037, 221.009225098777, 222.427421905688, 
    223.409043596671, 223.053118987031, 220.99400649008, 218.700089383387, 
    216.749433283216, 214.781942597731, 212.93733508912, 211.924255515429, 
    212.307635212884, 214.258016039856, 216.118916197104, 217.36439084234, 
    218.364655224643, 218.465958635915, 217.088890942368, 215.732558075318, 
    214.362379288544, 213.936827189486, 213.25196213963, 213.886884864576, 
    214.077968963099, 214.264940736677, 214.183193009767, 213.292519736471,
  210.874137236061, 211.12702694795, 212.32788195992, 212.655286375851, 
    212.846170771129, 216.165770783396, 219.700832829119, 220.211123807579, 
    218.343948264978, 216.543762131395, 216.068992292437, 216.857671810473, 
    216.577018152187, 214.107279054091, 214.659180773222, 216.497871269176, 
    220.441051659514, 220.332629136827, 219.801670643558, 217.85314885347, 
    216.566574518548, 215.432388137588, 214.48550854701, 213.543370765679, 
    212.480014117164, 212.12296771864, 213.757537621881, 214.802143150911, 
    214.006825180349, 215.764051056924, 218.639336478127, 218.917272328092, 
    219.622070364309, 220.452313389856, 220.765588959345, 222.053333979915, 
    223.076059845713, 220.729339982249, 217.11057883156, 214.881855217501, 
    214.423540712669, 213.587066094741, 212.214503234485, 212.691937574394, 
    215.095312783261, 216.995553690038, 217.334543190551, 217.32388177492, 
    218.063386515043, 219.403941753119, 218.253898231529, 216.727000680873, 
    213.831137460343, 212.774944058929, 211.741102634007, 210.189944146933, 
    211.676276465396, 213.799670751424, 213.933551331462, 212.562537487296,
  212.06082491118, 212.578671288042, 214.441414510291, 214.653872955708, 
    215.813250290574, 218.308120064011, 219.91088705548, 219.073978878691, 
    218.649647973651, 218.401465304764, 219.354572249207, 221.16112872008, 
    219.571448505749, 215.41152625416, 216.267109628988, 222.151184745685, 
    222.809029108404, 222.863497308812, 221.080287074623, 217.853357857546, 
    216.922943077993, 215.477235561819, 214.420535928838, 212.488789765495, 
    210.216684697294, 208.769604448671, 210.019201535634, 212.221435346268, 
    216.46365069443, 221.222675573765, 218.605826714776, 215.817550862907, 
    213.830597683851, 213.50558094528, 212.968428149748, 214.824349537775, 
    217.196150076553, 217.644354844307, 215.869558384757, 214.030802492706, 
    213.425390392558, 214.005369817386, 214.654547064063, 215.968267713553, 
    217.479632948083, 217.84627957648, 217.723779178364, 217.796112325405, 
    220.088567816102, 222.229539194377, 219.291097086639, 216.087966845463, 
    213.734511742776, 210.911179717645, 212.874574527187, 212.899273956693, 
    213.150663183803, 212.580921777469, 212.287938350387, 212.588544925405,
  216.862318900379, 215.898763784151, 215.892903086348, 217.302406391965, 
    217.972692692789, 217.7095398754, 219.653166668887, 220.807154972293, 
    220.026760596421, 219.581522256805, 220.950204279572, 223.776073105271, 
    224.270605467513, 221.795482612826, 215.617940881716, 219.218093585454, 
    224.308761939847, 223.231691415778, 219.604297478271, 217.934974648335, 
    218.523118346246, 217.5162528005, 216.898502342114, 215.832759074423, 
    213.447699010393, 211.888980800585, 212.494254642298, 215.546033393471, 
    220.468050929705, 220.982594582312, 217.770675649831, 215.187015501041, 
    211.720131426603, 211.909462752803, 214.351188087011, 216.704369514461, 
    219.67952955376, 220.587710441458, 218.881003787643, 216.923677600139, 
    215.321981804727, 214.799942899032, 215.215342708228, 216.534932506309, 
    217.378932760592, 216.654866171248, 215.887527466752, 215.944675228374, 
    216.626507099432, 216.014916471423, 218.745553746435, 220.966695600268, 
    218.837212188222, 215.194797879021, 213.827156479976, 218.631224770572, 
    221.390589518107, 221.185569944145, 219.678786116247, 218.274281149718,
  222.307521026736, 220.793030728109, 220.134019750161, 220.274455810409, 
    220.442113215891, 219.936598684817, 220.342776988656, 220.254931871867, 
    221.456118674438, 222.605026794218, 223.31201941323, 222.878714186416, 
    223.985658751365, 226.073822178039, 225.220209896662, 220.201364584374, 
    219.910604758514, 224.629102514918, 226.342805196552, 225.413353068712, 
    225.56844611703, 223.872054304125, 221.196388391708, 220.015089048294, 
    219.526324524554, 218.880922614212, 219.022231603404, 219.819082330239, 
    221.533059191261, 221.911084703746, 224.030756909912, 224.52292392534, 
    220.844375988075, 219.330737666608, 220.344336119826, 221.040572598062, 
    220.26890162628, 219.276300655844, 221.273846240605, 222.500571534569, 
    221.185821458339, 219.653064876042, 218.702256143919, 218.308164147263, 
    217.722179141084, 217.891790878432, 219.870260125152, 221.66547323859, 
    222.236078810557, 220.945778669185, 218.897830953082, 220.045161092487, 
    220.90276079089, 221.454620936124, 219.315911652661, 218.045342796818, 
    220.365650664613, 223.707342956961, 225.014129806996, 224.234615457835,
  225.368582068254, 223.199755669581, 221.101110217648, 221.808377528771, 
    223.717322842591, 223.329150984208, 223.578828294454, 222.881025398954, 
    221.687526379388, 222.657515483493, 224.51732116942, 223.865989627093, 
    223.790768373073, 224.679715968875, 226.786762243393, 226.371127961349, 
    221.244685180983, 222.31596377864, 226.333321613364, 229.221995622067, 
    230.586537991473, 230.552261136045, 227.665423117146, 224.784242199923, 
    222.56101051156, 221.698170146508, 224.73684605489, 226.240682275386, 
    225.388080501076, 225.355696651387, 224.245417346736, 222.941927734357, 
    225.369560286335, 227.806105806344, 227.74997795041, 226.814739855197, 
    225.109579331178, 222.322925783579, 221.372957676891, 222.341765048868, 
    223.829234730768, 224.269052604776, 223.046255429498, 221.558244998391, 
    221.57996487713, 223.201689667779, 225.221310394394, 226.4897259992, 
    227.431623484529, 226.656549511669, 223.643941435849, 222.552541518981, 
    223.329307537057, 223.567891314832, 223.276273832426, 221.456985798217, 
    219.727837771662, 221.761291219371, 223.48139082911, 225.488786293125,
  224.646309897674, 223.791914919594, 222.038954193276, 221.643414002942, 
    225.491517671811, 224.757842046067, 224.528252813008, 224.552973722145, 
    222.833802804669, 223.856491175604, 224.700899666732, 223.877953180274, 
    224.989635540188, 225.41613588171, 225.651666740002, 225.635662827234, 
    222.802450308507, 223.360628005806, 224.503446667155, 227.384383464741, 
    229.773616806221, 229.000124822283, 226.880686924024, 225.795648934923, 
    225.220137781502, 227.143486524089, 231.715446557335, 230.513269886061, 
    226.644917642181, 224.771082305911, 224.461500283668, 224.959764868137, 
    226.496318191256, 228.061204875991, 228.93970711412, 227.377327702455, 
    225.370857981567, 224.193300795737, 222.909054567166, 223.58674141281, 
    225.685208893567, 226.261665509597, 225.34624896687, 223.381063014255, 
    222.900041896624, 224.694964668123, 226.641462984073, 226.953719886692, 
    226.591510147088, 226.492989730658, 224.340109921364, 223.726043932358, 
    226.779020940453, 227.139774870799, 225.183896203544, 223.830839259339, 
    221.309041451345, 221.74098203823, 224.416328130366, 225.912703939132,
  224.129965079442, 223.545114234248, 221.66189594992, 221.812458223146, 
    224.482787410095, 224.124452415284, 224.003712482179, 222.932348249849, 
    221.961338110802, 223.235201447706, 223.489553676971, 224.242653593433, 
    224.239364775781, 224.398413388034, 223.71179534251, 222.608228683792, 
    223.746730906827, 220.069321653437, 224.106101028769, 226.64793361948, 
    225.949390191135, 224.174813837675, 222.667183808171, 222.764263892964, 
    222.808417908338, 227.515148192525, 230.79800050022, 228.22780747363, 
    225.138743850379, 223.050691429508, 222.505192069536, 222.60904499068, 
    224.658970779897, 226.333848265509, 226.678607114221, 225.310119604228, 
    223.406524554594, 223.05995802114, 222.864531457002, 225.05951088738, 
    225.733505082032, 224.74455188517, 223.474411580916, 222.394226031633, 
    221.755351697299, 224.572054818194, 225.549770374791, 225.968376141322, 
    225.713844495897, 225.127751910191, 224.157339706092, 223.552494311281, 
    227.171829688454, 227.523501374875, 224.393594612909, 223.730380802615, 
    221.871690827815, 221.117870030709, 225.528414285949, 225.85488371562,
  224.144762522314, 222.784435520363, 221.342551105727, 222.768252904108, 
    223.408261488668, 223.870497000439, 223.576706837815, 223.081372955454, 
    222.558662256698, 222.223980320981, 223.812385748302, 223.725176036488, 
    223.667304215322, 222.579128939381, 220.641113324087, 222.894790977239, 
    220.08656274693, 223.129808322471, 224.741971969717, 224.308883402895, 
    222.4698063058, 220.992023221399, 221.792729323237, 221.556843019748, 
    222.055724914399, 226.465820624159, 226.488856817604, 223.872099164854, 
    222.535686326902, 221.739470272122, 220.955721159898, 221.934531758614, 
    223.961498739945, 224.770969106778, 223.908430536907, 222.242812861118, 
    222.083579635557, 220.725428143884, 221.526217037568, 224.319477068207, 
    224.293931383154, 224.120704667347, 222.652733955114, 220.731102676266, 
    222.474285864763, 223.835778637902, 224.130241590312, 223.394020347393, 
    223.229693695251, 222.786747251515, 221.368206590071, 222.382741864528, 
    224.596865248423, 223.965364435926, 223.126708143878, 221.652804544362, 
    220.513923019621, 222.572782629203, 225.878559419711, 224.903796341488,
  224.854548884476, 224.234355355225, 224.062407859029, 224.639159960991, 
    225.121210280219, 226.435900841447, 226.766192700827, 226.353732837167, 
    225.847637894109, 226.412602113592, 225.964089453941, 225.459542287683, 
    226.291085725674, 224.4162633984, 223.268204722417, 222.438493685585, 
    222.519329912556, 227.187159053698, 225.18667855181, 224.505482469914, 
    225.582839178137, 223.293752145976, 223.409931517959, 222.522400492026, 
    224.837116330069, 226.55250802998, 225.338877394185, 224.851427777745, 
    225.859486337261, 225.568757307528, 224.975236394559, 225.530940312657, 
    225.445037666378, 223.631007935832, 224.407357265813, 225.662905645469, 
    224.269383359553, 224.283348462578, 224.206196075652, 226.014584797996, 
    226.666513612639, 224.666387981291, 225.13138270375, 226.125572014692, 
    226.553894490379, 225.847279351028, 224.948928086668, 225.304424169597, 
    226.000325758052, 224.870773520587, 224.655098304269, 225.32481386629, 
    225.779846710054, 225.197054754597, 225.61995280433, 224.870122885657, 
    224.246295022642, 225.254051886029, 226.02614135453, 224.879031439747,
  226.162698030489, 227.264618813215, 226.846839127549, 228.200619225618, 
    226.777492173459, 228.680612411229, 227.792361904258, 228.324887871608, 
    225.995446171695, 229.138200546685, 228.963792398187, 227.901968924991, 
    227.265075513305, 226.739396122048, 225.658470813962, 226.342540783014, 
    227.783822529747, 225.828204610379, 225.875767585661, 226.280909778206, 
    228.720561370488, 227.451001927973, 225.113397184642, 226.2923926023, 
    227.342924011941, 227.475799256991, 226.681862866363, 226.235524809201, 
    227.869016217702, 228.473705526116, 227.59281079449, 227.222949262954, 
    227.314402330801, 227.034155517005, 227.268198649982, 227.634874046276, 
    227.432383963346, 226.9746084652, 226.799923042635, 226.405467332688, 
    225.915677997245, 227.62742203395, 228.83351186752, 228.471346652126, 
    228.19151637841, 228.162388766734, 227.634249150042, 227.168072901254, 
    227.018977700299, 227.090586139963, 227.335523616728, 226.968048355221, 
    227.472077060242, 226.813120204723, 227.045325466488, 226.624392739256, 
    227.471425717503, 226.351057000273, 226.983372565539, 226.210202326877,
  225.614020661528, 226.639016292852, 227.773515217286, 227.693179563281, 
    228.665816305609, 229.307364281378, 228.83742986919, 227.738522311278, 
    229.95872869171, 228.523261839303, 227.671470798456, 227.867004093239, 
    228.115431654752, 228.169072446751, 228.104869349064, 227.749076550632, 
    228.682525451925, 226.85844681338, 225.707225801928, 226.679729002168, 
    226.172176230786, 227.502355230151, 226.908546519605, 226.823453538074, 
    227.517704729485, 226.876847315668, 226.249835140541, 227.185427194257, 
    225.96445538092, 226.178695991015, 226.326122353179, 226.708209097842, 
    227.106438505271, 227.643549896744, 227.451947081001, 227.536797633374, 
    227.367112126434, 226.957765534618, 226.74943245774, 227.060601789017, 
    226.905660511132, 227.538575989803, 227.527021769, 226.389663427538, 
    226.235154156485, 226.752096909267, 226.900204901372, 226.970129912726, 
    226.964487295928, 226.904758067761, 226.8596235797, 228.485696622735, 
    227.570255181424, 226.48904448293, 226.555036916015, 227.221819620198, 
    227.382629922156, 225.837006678393, 226.920598642331, 227.117028910489,
  227.106301844462, 227.824566080852, 226.778094107016, 226.634519228788, 
    226.94789234971, 225.927576773456, 225.368548850498, 224.767681962329, 
    224.118038988306, 224.354554052257, 227.586668248593, 227.096170445178, 
    226.797276527415, 226.935140572718, 226.691365743786, 226.484914519902, 
    226.364163866639, 226.268850671789, 227.46864763122, 227.033375521263, 
    226.722236896471, 226.299073838001, 227.401685867888, 226.467995172367, 
    227.059710998291, 227.005126786187, 226.309604976006, 226.766191052841, 
    225.795125669633, 226.651228540262, 226.544481731119, 226.042160513202, 
    227.547138093592, 227.958716322737, 227.904414090707, 227.78117527157, 
    227.480910511528, 226.911086875106, 225.855350189291, 225.695167957178, 
    226.618732199403, 226.845780188258, 226.090796601953, 226.143298339078, 
    226.891910541925, 227.534603431797, 226.950021340244, 227.245885184487, 
    227.55900756878, 226.256280086407, 225.862716182158, 227.922794370754, 
    227.911238572307, 226.865614340654, 226.5869458166, 226.251633518066, 
    226.325381856748, 226.472528121257, 224.198771829211, 225.494239709554,
  232.021341577941, 228.547444947743, 226.825415191698, 227.380066224059, 
    228.57695932619, 227.027135471747, 226.710342441116, 228.031838962848, 
    226.459991744526, 225.755056865725, 225.398506948606, 225.667376562534, 
    227.189646386019, 227.447146723813, 226.716214581965, 226.519186204017, 
    226.533990042982, 226.796738829815, 227.415643198236, 226.608428401247, 
    226.657943972742, 227.193007213699, 227.46857510821, 227.079157349173, 
    226.940337101062, 227.374521231879, 227.317207537236, 226.12954870648, 
    225.466250259186, 226.308377103059, 227.796975811172, 227.866288847489, 
    227.007992674201, 227.262463214728, 227.462845877457, 227.836129280888, 
    228.331007528917, 228.103206779401, 227.175770150064, 226.85551349871, 
    226.490256394442, 226.245199954622, 226.653024538228, 226.413541687225, 
    226.657244438128, 226.741574909763, 226.814531536848, 226.869485018288, 
    226.651151373008, 226.907188713106, 226.780999538501, 226.959106635639, 
    226.740727570242, 227.092383472693, 226.537521665511, 226.833446446603, 
    227.025704263093, 227.060965901046, 226.07670663147, 223.94577633116,
  224.97821540615, 224.466917270858, 225.440029651145, 225.773526963094, 
    227.039855096594, 227.012708945747, 226.347208046774, 225.159820486113, 
    225.406453250534, 226.150563237193, 226.310260148522, 225.02998242731, 
    225.10931057803, 226.829618550568, 226.552975099033, 225.881800625464, 
    225.479250527565, 225.282054392818, 225.947214076487, 226.025233879078, 
    225.308257554347, 224.578259229056, 225.079357354832, 226.317998682399, 
    226.799957278804, 226.15359067308, 225.544950194252, 225.715171895329, 
    225.068286970704, 224.472741209349, 223.22834052624, 226.370354656952, 
    226.835826749688, 226.176481440718, 226.224515397423, 226.219493542058, 
    225.722751672493, 225.507347911612, 225.596597004384, 226.383872666667, 
    226.02907508023, 226.026853064197, 226.194885936396, 225.861674047549, 
    224.730511688905, 224.081296575916, 224.733250500371, 225.616255128698, 
    225.444273577576, 225.544939160164, 225.849360412462, 226.057313938771, 
    226.243788242561, 226.622559394562, 226.637111035637, 226.179645873401, 
    225.14580442551, 225.137242476773, 225.666318849303, 223.395480309745,
  222.750249799365, 219.77117657562, 220.916568083833, 222.810766574327, 
    222.884000030683, 223.387546247677, 223.687780006286, 222.382982150242, 
    221.402974138619, 224.603362087963, 225.274491813565, 223.980973052481, 
    221.378776490988, 221.98743528189, 224.316424025744, 224.555199338034, 
    223.625775146422, 221.470606275183, 222.397429017513, 223.763750537704, 
    223.565766410203, 222.470514287516, 221.19261296892, 222.542864240638, 
    223.543393859915, 224.235083386307, 223.763167527128, 223.146721805043, 
    222.552344154705, 222.954853782555, 222.697196241242, 223.200229366282, 
    225.122147029306, 224.522526898276, 222.918621011411, 222.233450989393, 
    221.326693807794, 220.306219516416, 221.310307170463, 224.171707913418, 
    225.723556554418, 224.597308373136, 223.010104585142, 222.783204461393, 
    222.89853922196, 221.927680213218, 222.306665502096, 224.363150293095, 
    223.58647562898, 222.913790769879, 223.53953718295, 222.497029597748, 
    221.730765302945, 221.960568973236, 222.144339000269, 221.795519001719, 
    221.039259687512, 224.762671718422, 224.388735555843, 223.272882360825,
  223.061549823793, 222.472931852855, 222.226507476758, 224.608967037773, 
    223.446004060688, 222.185524825669, 221.938405943875, 219.614248368186, 
    217.889863759681, 221.929723797124, 226.247379533299, 224.483670142878, 
    222.539334172601, 220.632545071227, 220.881688274145, 222.233431665128, 
    223.200162624338, 223.526606315377, 222.33085771064, 222.487128815005, 
    221.137590627099, 220.206797882761, 222.866901420834, 224.410249598399, 
    222.06939978261, 220.377508170663, 221.435589582296, 221.896293059063, 
    222.354885576497, 222.514968482318, 222.587250054726, 222.919875949465, 
    226.02015810014, 226.103048978713, 223.533549534683, 221.023411422173, 
    219.433460678994, 218.473032925701, 220.319720652535, 223.761338295462, 
    226.532190301777, 225.546465112525, 223.83973114291, 222.250165616749, 
    221.707451906676, 221.528626982591, 219.544983098463, 221.860021260609, 
    223.843732220476, 222.935036812825, 223.408691367301, 223.951118970386, 
    222.538951799199, 220.790287950297, 220.517245985067, 219.394044539517, 
    220.22290232035, 222.930739136459, 225.960688684598, 224.640447448985,
  225.051167610955, 224.389344461712, 223.843962936705, 226.243183227111, 
    226.094957227896, 223.785161554485, 221.607285249641, 220.03435452257, 
    220.404296890415, 223.481162163623, 228.518871334336, 227.978186121108, 
    224.011890585157, 222.536858362559, 220.358964333087, 219.384267019847, 
    222.761553122332, 225.007822253986, 224.722442898973, 223.300225694287, 
    222.363077861006, 220.669678242272, 221.646813010022, 225.789373480822, 
    224.918455543977, 223.615699062774, 223.22093005106, 222.261758830128, 
    222.054652497641, 222.219772491098, 221.5043923829, 221.166769345131, 
    224.673818890086, 228.278903976072, 227.19755273702, 223.907232565715, 
    222.503172137013, 221.494933980005, 221.825036658842, 224.52512595955, 
    226.994848213622, 227.679964951996, 227.022528220083, 225.216117000827, 
    223.981733121172, 222.478831246455, 221.763535886298, 221.938967601555, 
    224.055529053789, 223.512998893704, 223.934307471292, 225.59844116006, 
    225.06907231967, 223.691964448393, 223.074939382359, 222.592692967118, 
    223.528034454466, 225.49012047088, 227.435549256154, 226.271636632971,
  222.299654424769, 223.097643327346, 223.123719291122, 225.623425319152, 
    229.642461186599, 228.081323915144, 225.61759213694, 223.690134155175, 
    221.681537705457, 223.292027403546, 227.255595612929, 227.591861243428, 
    224.137917839081, 222.089730106729, 219.816805053677, 219.467872153364, 
    221.577000292649, 223.765725340983, 223.800128585894, 223.009221911196, 
    222.893117375321, 220.647705241207, 221.799460398895, 225.513354001626, 
    226.201039987441, 226.716738063247, 223.869150880337, 221.880989921339, 
    221.486150035921, 220.076743535595, 219.61017466421, 221.199425645945, 
    224.336132014113, 228.444074938285, 228.616224430655, 226.392987995245, 
    223.546766419529, 220.870814569549, 222.067059364135, 223.818811773071, 
    225.992311900546, 227.361051012175, 226.968177976445, 225.716080063272, 
    224.269699026567, 221.77302586577, 221.46072514427, 222.499648614493, 
    222.853720916667, 223.443657569868, 224.845746069291, 225.969454544621, 
    227.580715917303, 227.070398844552, 225.38103164929, 225.163771770309, 
    223.837192058352, 221.704206260414, 221.94986850471, 221.867602408963,
  223.853062477399, 225.631295842449, 223.922906350355, 224.950644513319, 
    226.336061699581, 225.625234100443, 223.296428258642, 220.207484035721, 
    220.623208008288, 222.7942890383, 224.426066348518, 223.90818582531, 
    222.194685887892, 220.478654906254, 218.834716314582, 218.324247753777, 
    219.212510145105, 219.840409534683, 220.23231917806, 221.269675411332, 
    219.793858274808, 219.501461208007, 222.150497184893, 225.764257745012, 
    227.98201748224, 225.043583967074, 220.362244435825, 219.125026063372, 
    217.443942161228, 217.241284895607, 218.274966021452, 219.81137612654, 
    221.828339114932, 224.171816419172, 224.193705011534, 222.960631976737, 
    220.566777632296, 219.770643464684, 222.345359243997, 223.205265357718, 
    222.784603699855, 223.18307211236, 223.732935652758, 223.446213266219, 
    220.919493395338, 219.114916876097, 219.266977215717, 220.78802798417, 
    222.461592362272, 224.201488965508, 226.425003498744, 227.491572007954, 
    229.376513083172, 230.363036684341, 228.277479292323, 223.828867908021, 
    218.989272325335, 216.801368901277, 219.361237445303, 219.366868535478,
  218.388399759949, 217.46014951134, 216.889516265531, 218.080789350392, 
    219.063610185158, 218.821869930088, 217.07877160561, 220.988402055738, 
    222.375390300796, 219.910656407411, 219.340145460363, 218.808136676046, 
    217.749667983355, 216.65523072287, 216.461517657111, 216.630656954255, 
    217.81083371355, 219.356708849524, 219.567483921084, 217.973592059478, 
    220.435068469453, 226.68738636393, 224.360764039381, 220.071140358253, 
    220.052706567413, 218.449275162857, 218.554691847876, 217.679785201144, 
    216.293456281067, 216.920294939066, 215.773039338807, 215.207073552452, 
    216.320200231093, 217.41184071003, 217.559710664534, 217.317224260719, 
    218.494800157599, 220.640383600346, 222.150348123614, 221.343206790348, 
    219.717819616619, 219.796096067723, 219.724628125953, 218.143054425572, 
    216.696451899573, 217.554081258882, 219.084003140489, 222.073311322315, 
    219.164787929581, 216.395451162838, 219.46436641897, 220.1358203628, 
    221.33976032305, 222.110681958446, 220.774820896403, 218.429794428702, 
    216.31681653339, 215.818637643885, 215.937660732124, 217.938610064675,
  217.052251459006, 214.368328280008, 213.207181957455, 214.858444203455, 
    215.445855387569, 215.066322656454, 215.693396294236, 216.125562767142, 
    216.464788546482, 215.280645760083, 214.615145277462, 213.994642016588, 
    213.531254570443, 213.873181915469, 214.515253797756, 216.204581182985, 
    218.424148550985, 220.505540803908, 220.529661640048, 219.391082586432, 
    219.115401728905, 219.191132664638, 217.852314573088, 216.811000719166, 
    216.984103778072, 217.145186623135, 216.351330837701, 215.257859377454, 
    215.60758802353, 215.849731020099, 215.172610126061, 213.690815274175, 
    211.761527317013, 210.301141605868, 211.302907851857, 213.510322225173, 
    216.042985558784, 219.998349236271, 222.551966762886, 223.798463802886, 
    221.054712503392, 218.040358205959, 216.393445654391, 215.111045934698, 
    216.720646461811, 218.162621306755, 217.308972514165, 214.069584752723, 
    212.027526609747, 210.441023545628, 214.405549900734, 216.372691824678, 
    216.735921490868, 216.878269313285, 217.924823031829, 218.784156249639, 
    217.521355136628, 215.484587781418, 214.717407050212, 215.4213967015,
  214.27528789683, 212.554079198448, 211.984867367751, 212.358945935338, 
    212.727081674569, 212.640750234626, 213.360047149822, 215.039629009893, 
    215.565606619546, 214.322735951193, 212.736928565703, 211.685076399891, 
    211.772763989297, 212.300487713465, 212.988134563062, 214.37576021394, 
    216.497172638431, 218.609920299102, 219.274877247666, 218.054278282275, 
    217.482695334012, 216.442333600938, 215.598926189677, 215.737330241034, 
    215.157356200193, 213.944573492066, 213.305435543145, 213.503918498479, 
    213.936502929779, 214.339537326897, 214.757461579991, 214.792540842484, 
    213.687532730245, 213.808266182969, 214.171413850363, 213.664803640159, 
    214.951298368603, 218.109209240877, 217.375018050801, 216.783458062113, 
    215.623277813983, 212.456498351983, 210.111434312994, 209.659925126478, 
    209.656454921039, 211.253820020532, 213.693826183076, 215.087529186924, 
    213.72979532919, 213.144780606994, 212.324141526617, 213.952483028885, 
    216.13634300715, 218.144519672365, 218.773231737146, 218.164657867066, 
    217.464647387259, 216.741908565906, 217.289634165886, 215.75283880757,
  217.108545959494, 215.680041006396, 214.374746788796, 213.487008050511, 
    212.874076771489, 212.867644306686, 214.210210792805, 216.053793711774, 
    217.293943926539, 217.093762025623, 216.258408098993, 215.251740211248, 
    213.964592147403, 212.963190058252, 212.449296800412, 212.727166233952, 
    212.711054372704, 212.420555738733, 213.335135881459, 213.973634764112, 
    214.058081298878, 213.972928446567, 213.895328448722, 213.075483983598, 
    211.562468910811, 209.922760514089, 209.043286909014, 209.372097172196, 
    210.66925729526, 212.40769974198, 213.754291831082, 214.695058087982, 
    215.589589960488, 215.498291029964, 214.637117431399, 214.276512603443, 
    214.937254942589, 216.682531130742, 218.244155336158, 216.812099968197, 
    215.3935205953, 213.075383236096, 211.417478207761, 210.09951606764, 
    209.049760070584, 208.867333065662, 209.221015090328, 210.921359676435, 
    213.479464887791, 214.012245884062, 214.091044965323, 215.043618622781, 
    215.401878457358, 215.906378440779, 216.501344331456, 216.744178119751, 
    217.629053499272, 218.568696672809, 218.901394959892, 218.464979038061,
  217.361929543541, 217.188381875635, 216.919812574403, 216.584133886829, 
    216.308643816665, 216.143718732867, 216.006663856848, 216.394023401209, 
    217.473177595397, 218.567713784539, 218.714228906038, 218.164554808722, 
    217.669206093231, 217.412111784595, 217.723490353716, 217.817765974013, 
    217.660423435814, 216.680592112431, 215.705577571772, 214.759705631447, 
    214.05940380486, 213.396351098719, 212.664295762936, 211.881698549593, 
    211.200956119826, 210.582168946054, 210.300036459584, 210.608617238564, 
    210.925349869415, 211.531202049347, 213.258164992344, 215.156969914901, 
    215.91666455334, 215.684718458216, 214.957920697186, 214.340083259573, 
    213.758909066057, 213.204973552483, 213.644786950255, 215.070093069661, 
    216.003250744411, 216.070627249334, 215.82836789859, 215.662145275837, 
    216.082134762379, 217.046877624366, 217.771592732944, 218.178441014936, 
    218.298707169834, 218.116034012029, 217.906101481231, 216.966935125036, 
    215.594514872721, 214.287212502469, 213.449303485495, 213.660491736538, 
    214.264160101457, 215.065613881067, 216.250320459482, 217.077675516553,
  215.060016558455, 215.512144314359, 215.611682722925, 215.539216021735, 
    215.462165488934, 215.434864392638, 215.665231861808, 215.914498387591, 
    215.906973843605, 215.812537325851, 215.869263394441, 216.002737572756, 
    216.037054099332, 215.944837232787, 215.733106666955, 215.298419425203, 
    215.182798510164, 215.252967904746, 215.186763784288, 215.203003067419, 
    215.137753352136, 215.003233108688, 214.948545131847, 214.829981871901, 
    214.703748458573, 214.793887552243, 214.740185806327, 214.609417300125, 
    214.800686840865, 215.343792230578, 215.569596512349, 215.416222001325, 
    215.307452206676, 215.185944369979, 214.913386880912, 214.533767133004, 
    214.252495416729, 214.114286786049, 214.342425244698, 215.106053967154, 
    215.895057697995, 216.529563982183, 217.031779395583, 217.442300553074, 
    217.73067720053, 217.671416421759, 217.491540527461, 217.424366978941, 
    217.601056004472, 217.768762248742, 217.579625112267, 217.164336283197, 
    216.695923843414, 216.175167726128, 215.874639766294, 215.655754597722, 
    215.027767904844, 214.268727308549, 214.078948251096, 214.486664491637,
  212.423374691385, 211.772527543186, 211.381178793962, 211.218076281596, 
    211.269394475872, 211.379787199721, 211.291103890016, 211.079447802615, 
    210.955824986941, 210.925461870953, 210.96087474643, 211.017337154342, 
    211.086478890729, 211.209371156175, 211.376624212215, 211.674415044856, 
    211.979214146487, 212.187785509386, 212.41200912825, 212.476140421509, 
    212.522994262897, 212.551566105984, 212.609004839674, 212.706838375976, 
    212.894209710255, 213.004822717318, 213.137439335139, 213.4141729513, 
    213.888904499848, 214.259995163397, 214.335353048548, 213.823856919323, 
    212.772582479241, 211.573755509041, 210.626316918957, 210.077832812003, 
    209.855129342334, 209.964375397336, 210.303544643213, 210.677342208585, 
    211.185724948698, 211.791073995809, 212.275814792923, 212.595861610591, 
    212.841704765587, 213.158623743836, 213.501611498802, 213.738500469551, 
    213.782759336879, 213.668090204165, 213.401661879005, 213.161688352517, 
    213.010554398095, 212.936125539511, 212.90045026672, 213.050355909262, 
    213.255638625896, 213.595073125632, 213.77208600817, 213.235831776297,
  225.568757939197, 225.799280680904, 225.888280151834, 225.736881096607, 
    225.429238530589, 225.05818968341, 224.788295689113, 224.657165637095, 
    224.808815144682, 225.132512252012, 225.508010391478, 225.767942986023, 
    225.952565289663, 226.056063148143, 226.079873109919, 226.051709283885, 
    226.061732371295, 225.957678110428, 225.800366296355, 225.828033463959, 
    225.834148832929, 225.879984154516, 225.9147263809, 226.156118618351, 
    226.548967616919, 226.764883688565, 226.653604579708, 226.584783512363, 
    226.795851639303, 227.164625931626, 227.526755901481, 227.621376965173, 
    227.32381679298, 226.809810230188, 226.329897152094, 225.904905393816, 
    225.61285271085, 225.442215751321, 225.419727045649, 225.461921347715, 
    225.594857898893, 225.75538147727, 225.911191232275, 225.968063952594, 
    225.933398075708, 225.896903829673, 225.858711333462, 225.730186717707, 
    225.524565159534, 225.27732411179, 225.042361899474, 224.921132554322, 
    224.87195734107, 224.863243334667, 224.874531534632, 224.891676475735, 
    224.948513641501, 225.033003600676, 225.158845099829, 225.330515166018,
  232.665914706398, 233.160035759717, 233.441491403379, 233.533184069146, 
    233.437659409465, 232.972343755982, 232.278573185223, 232.027359563793, 
    231.799635371797, 231.370690253624, 230.794027653735, 230.146035395345, 
    229.518633380424, 228.879231176, 228.250515251925, 227.62678039811, 
    227.206763990496, 226.9399309508, 226.947146494405, 226.764172987365, 
    226.491075950032, 226.290844156342, 226.17765304823, 225.940763607117, 
    225.114827820554, 224.196130900503, 223.914643517459, 224.184352535301, 
    224.872522760338, 225.32635180902, 225.57497081467, 226.004980099414, 
    226.266386250472, 226.296044546777, 226.453965672179, 226.900465409596, 
    227.470876771224, 228.157209570633, 228.855749489675, 229.332760469704, 
    229.324202271617, 229.123283654104, 229.482281708044, 230.403360972785, 
    230.269117001554, 228.908870152665, 228.003606595063, 228.047053639281, 
    228.27307775023, 228.358244413984, 228.43300583437, 228.611130727501, 
    228.89347627063, 229.186275346899, 229.445041906742, 229.875101928046, 
    230.261525652758, 230.649874689518, 231.259604234841, 232.023305078121,
  233.534017157154, 234.47427840045, 234.577470818424, 234.100464147403, 
    233.409430606025, 233.162174872873, 232.945452653393, 232.250080679644, 
    231.983024661795, 232.242429877547, 232.692843078363, 232.857187232467, 
    232.930645276173, 232.59120812598, 231.832565780279, 230.790205717985, 
    230.082178439046, 229.463792040564, 229.610216061278, 230.017841819944, 
    230.351775144736, 230.564697825471, 230.552811188665, 230.111358357132, 
    229.356936744931, 228.909142361678, 227.816279865668, 226.904184285494, 
    226.29245549138, 225.977974922303, 225.871025209754, 226.245330076085, 
    226.702757381213, 226.963902734359, 227.548517738141, 228.439307668171, 
    229.312044334626, 230.141584479027, 230.995418274678, 231.938087794132, 
    233.016939556499, 233.957627499851, 234.122817769985, 233.950262896385, 
    234.19794828018, 233.414857244032, 231.411239709592, 229.770405935077, 
    228.911937519023, 228.94311894251, 229.612348851367, 230.809889737461, 
    232.161203222087, 232.489532409995, 231.711340470181, 230.750026807269, 
    230.697119688503, 231.154414193416, 231.690006038443, 232.448160043084,
  238.255898323034, 237.392574646292, 236.41899679487, 234.382012144933, 
    231.711940559829, 230.650493037288, 231.820406483415, 233.064917489616, 
    235.039529165309, 237.215007365291, 239.538655902591, 241.171032357576, 
    241.390071424071, 241.825329923802, 239.914070711587, 237.57388683448, 
    235.459132707808, 235.109994195389, 235.998912120912, 237.254556381422, 
    237.623202611073, 238.016057050035, 237.820883610367, 237.325826747314, 
    236.738998569857, 235.103378572403, 234.183670172395, 232.193691446152, 
    230.755427557667, 232.139169713818, 232.295387206392, 230.706816807952, 
    229.670409209728, 229.135639655853, 229.126584916031, 229.629278350815, 
    230.353512376309, 231.858503731923, 233.627831605206, 234.865216576101, 
    236.111356496956, 237.613133704453, 238.579465850092, 238.261899999852, 
    236.883340107543, 234.619565930378, 232.644013655319, 231.360687420421, 
    230.700690846647, 231.81067796287, 234.829727995096, 236.476068206796, 
    238.368225467124, 238.675525633143, 239.814379585168, 239.258633388024, 
    238.911972726671, 238.780832165848, 238.676555517983, 238.649261803866,
  241.92449140618, 240.971654366108, 239.259566356267, 239.415567116201, 
    238.470365704223, 235.51797758839, 234.64083839964, 236.194256640597, 
    239.96996642263, 244.587732360147, 247.234970869478, 245.789602849463, 
    245.226644784287, 247.239715144591, 243.893122353465, 239.781594187689, 
    237.875498618682, 238.850468139533, 240.176471656895, 241.810903792178, 
    241.81249589264, 241.689346885164, 241.345722202819, 240.966678114413, 
    241.484775377471, 240.854801481622, 238.620107113126, 237.76404042209, 
    237.493826772526, 235.434334370145, 234.687016909768, 235.630885729715, 
    235.465537591557, 234.399890183205, 233.726210182378, 232.609753283611, 
    232.472644276832, 234.821907865919, 238.790028002572, 240.986267705841, 
    240.878483976025, 240.323185024481, 239.896369116727, 238.129333222648, 
    235.581098042805, 234.367428222559, 235.262263468759, 236.314832945767, 
    237.012141661547, 237.383953125501, 240.052987306276, 241.244817411514, 
    243.474363530424, 242.45545261804, 240.896373786052, 244.396235957132, 
    243.802635025692, 241.174743381566, 240.673777752244, 241.195829898107,
  240.82316091579, 239.937308207433, 238.705948762509, 238.060123151753, 
    236.852352254582, 235.342734052197, 234.980797645678, 238.483635060699, 
    241.767392740785, 244.96590241856, 245.663462110338, 242.907894594066, 
    244.503686736214, 247.479400812395, 242.989224671673, 238.467608320438, 
    236.964162401655, 237.854403569579, 239.838353554446, 244.087445478271, 
    243.935651274341, 242.883749453692, 240.8091704331, 241.433015931307, 
    242.678304794962, 243.492884900438, 241.702931565495, 240.224418645255, 
    237.848055504049, 234.616202348269, 238.963059872307, 243.100145696983, 
    244.020212648034, 243.682603495378, 243.304771605426, 240.079291669643, 
    238.540158175358, 239.957953216458, 241.549065000604, 242.491810478956, 
    241.886858979115, 240.274074363739, 239.204167053757, 237.93494261915, 
    237.008059679312, 237.669531718428, 238.524815290499, 238.857287656117, 
    236.583290915913, 235.71063832166, 239.644131129092, 241.532127689443, 
    243.263543125492, 244.328486734432, 242.380334863256, 242.846451721044, 
    244.14286769503, 243.897292462492, 241.947835316181, 240.847819044025,
  241.736647899063, 241.258069082494, 240.609921342749, 239.451335455984, 
    239.270534015898, 240.181383470193, 237.604902263411, 237.320710397366, 
    240.21616831739, 243.601320461807, 245.196666548054, 243.14111564131, 
    241.90773609013, 244.816279077051, 247.943627553403, 242.06313088085, 
    237.62010200015, 238.115917180004, 245.30459296072, 249.281498113148, 
    247.244611394985, 245.870062941714, 242.658326249002, 240.79319102879, 
    240.656603331306, 241.674902935691, 240.790303861688, 239.291615885683, 
    237.372951828765, 237.910171292274, 244.70625749001, 247.151949016911, 
    247.591822494778, 244.284576670462, 242.602288475904, 240.79414216715, 
    240.127705311712, 240.448803287784, 241.769026292427, 243.219404111003, 
    243.429888530332, 242.438445735926, 241.285957638535, 239.935571625033, 
    239.732746821631, 241.61722382585, 243.945077805055, 245.091980736723, 
    245.002243175294, 245.505634273126, 242.341864687139, 240.462633082768, 
    242.785312976253, 244.166109700962, 243.222410929481, 240.204843277701, 
    238.31717238215, 239.234619118614, 242.174873109714, 241.871910325332,
  244.445311433742, 244.79370003234, 244.255002636057, 242.70520441546, 
    242.710047471943, 242.982185017912, 242.319379223935, 243.085918600648, 
    242.987000166071, 243.98787823893, 244.755522067346, 245.11762950759, 
    245.128026340095, 243.540699530721, 245.538357882128, 249.367372571169, 
    245.655849881062, 241.751754532406, 241.546625463279, 245.433187437224, 
    247.288765917749, 248.183640252281, 247.28102299727, 244.398615006782, 
    242.396942183255, 242.068297944161, 241.996353084952, 243.158906204149, 
    244.042512859085, 245.717076549301, 242.061423125938, 240.968549790577, 
    245.808522127, 245.454208845109, 245.06465890597, 244.957527016008, 
    246.779828146116, 247.901668668186, 243.560134936779, 241.629925556568, 
    243.330685130372, 244.720673389218, 245.022193982526, 244.859669325389, 
    245.77419927318, 246.874332419116, 246.629206826059, 246.092781979309, 
    245.797322031443, 247.555450092358, 248.009951958792, 246.909392035717, 
    245.420767790903, 244.59289722648, 246.651155439226, 245.649837537716, 
    242.977064318604, 240.521685574003, 239.985850314373, 242.512366348467,
  246.228562269257, 248.295105596421, 249.948607996427, 247.381748117297, 
    244.953104037636, 245.734071322408, 246.220010002711, 248.846997687793, 
    248.51338046688, 247.531900343907, 247.981773862238, 248.209948412954, 
    247.638452920307, 248.993095543789, 247.661362567881, 249.110518682962, 
    251.054072289192, 246.770255773011, 244.668739558426, 245.245004258403, 
    247.388983718775, 247.909290521665, 247.283046924793, 246.852965258395, 
    246.790847924977, 246.872284354913, 244.684130538756, 246.140220880729, 
    247.964116813996, 247.486151006297, 248.208816017165, 249.549709586263, 
    246.441012233134, 244.600909965031, 245.218244472837, 246.865949556007, 
    248.33435403657, 250.23255154289, 249.427547142158, 247.035196253054, 
    245.575761683868, 246.279476001548, 248.252826828405, 249.057033951403, 
    248.451236676236, 247.786486723233, 247.484425750742, 247.660515101218, 
    246.348443922833, 246.232521804168, 248.895677096705, 249.155935382623, 
    248.396283251128, 248.389129522352, 250.432071052822, 252.399228385461, 
    250.33155810376, 247.023362404738, 245.513705176029, 245.715679134132,
  251.141354312338, 253.681170644083, 254.298211736284, 252.09772453634, 
    249.92269651184, 250.338529269943, 250.423293591258, 251.815757970628, 
    252.577479363533, 250.149730611696, 251.112545759301, 250.622479595245, 
    249.458314333364, 252.611327413362, 251.713264665471, 252.15588065856, 
    253.410289241272, 252.622186688004, 250.317302263419, 247.57077897669, 
    249.215692266502, 251.146072314752, 251.237992558428, 251.908182232651, 
    248.449970409179, 244.899129916536, 245.171817040487, 249.374612629629, 
    252.503015833934, 254.540820806651, 254.069289770025, 251.822031015271, 
    250.567203083744, 249.041443460691, 248.603955087998, 251.422729161155, 
    253.027847550086, 253.184487563905, 252.280224447621, 250.522692145757, 
    249.830574279676, 250.05893364355, 251.76899021432, 252.816714237227, 
    251.544736501728, 250.224454975806, 249.658060043506, 249.239401629224, 
    251.049320731635, 252.036582117998, 254.535596203835, 253.157621935321, 
    249.360720998689, 252.164699627209, 254.245167133624, 255.076769283418, 
    255.991763748838, 252.381746107441, 249.333697117048, 249.339319970966,
  255.956005522941, 257.029343592463, 257.257493065667, 256.448347163506, 
    255.038253759196, 255.222153726819, 255.712812864528, 256.718531567844, 
    257.038463682356, 254.835577886362, 255.467744213259, 254.871575136247, 
    254.816282353659, 257.103348445972, 257.503914556491, 256.238186013092, 
    258.240832653159, 257.403153790008, 254.53503607539, 254.142650057208, 
    255.887772524339, 258.355282139563, 257.885520683479, 259.029338972974, 
    255.761947374394, 252.057262652524, 252.122355803079, 255.955982845801, 
    257.989032233592, 257.922560751741, 258.182647608013, 257.157979762276, 
    253.688152018401, 253.343299565579, 253.891671391741, 255.011231892216, 
    257.065611816671, 256.182028675136, 256.162299151154, 255.241864640828, 
    255.08931933027, 255.428685301157, 256.774972767294, 257.466657638417, 
    256.734426434984, 255.20324739746, 254.999814035519, 254.189801487326, 
    255.621707374637, 256.035767363431, 256.261741564642, 256.876199061308, 
    255.851342499988, 256.245118338468, 258.800008662789, 257.914988784147, 
    258.825275803725, 256.621326113463, 254.446109994154, 254.878203399383,
  257.648087927787, 258.690748841093, 257.312498202296, 256.912539697713, 
    257.245390766893, 257.118465389165, 259.22224989604, 258.12806089029, 
    259.400175716622, 260.290900584393, 259.124204685781, 258.930736480644, 
    259.320977038562, 261.360261298524, 260.294308956838, 258.441237187033, 
    259.709126867518, 258.118962988083, 258.869259211189, 259.091865433352, 
    259.503431402639, 260.795987639491, 257.901926554568, 259.625983506356, 
    258.560268059245, 258.650824309513, 257.521441782169, 259.710273189469, 
    259.465727432165, 259.748078941884, 258.284634360576, 257.184908459607, 
    256.265240149997, 257.455293260058, 257.558725400194, 257.646435507833, 
    260.658715718542, 258.797509604383, 256.250756457593, 256.082051377308, 
    257.349077864249, 257.093752919692, 259.114497181035, 257.63148606794, 
    256.835492834546, 257.092260043474, 258.335436252242, 257.279724647177, 
    258.219295822734, 260.153775766417, 257.916978607102, 258.843272550973, 
    259.471659677153, 258.383559111848, 260.377657344411, 259.306972984401, 
    257.595109339761, 257.456095524599, 256.590261561971, 257.653865224016,
  258.647584276629, 257.96784531896, 258.055597691628, 257.600197747934, 
    258.204147247377, 258.062782042482, 258.978340804994, 259.428803703621, 
    257.696483111642, 259.129960820958, 260.026727473926, 259.03738414906, 
    257.73890186144, 259.828051616702, 260.51079832333, 257.991980303716, 
    258.946950481505, 256.634793346681, 261.210192270301, 257.604674741234, 
    256.085303673155, 260.28394790032, 258.712866491664, 258.347709235995, 
    259.369656231606, 259.485578800831, 259.087094497206, 257.555855049803, 
    255.608382922744, 255.996851870588, 257.289448875058, 258.045008399194, 
    259.628286868436, 260.113006931194, 257.052593553808, 255.520502366252, 
    257.440262860713, 257.417147560487, 257.872678260279, 256.658788792516, 
    257.515921570424, 258.015273482141, 255.808718171991, 256.660683846066, 
    257.30587325751, 258.487007667164, 258.54330581859, 258.268743621395, 
    257.723264783169, 257.788843848666, 257.203389713531, 258.923731038756, 
    259.001704463116, 258.952084341709, 257.2051611026, 258.087423218108, 
    257.229616341214, 258.182253139486, 257.633821147032, 259.512000496773,
  259.031843451435, 257.954081623442, 258.056180906717, 257.449320595673, 
    259.52536389775, 257.844197740047, 259.455031519008, 259.384391347698, 
    260.688051806052, 256.734055973434, 257.904108129136, 259.378538606745, 
    258.429991254438, 258.440137014501, 259.429305974471, 258.075870943859, 
    258.586291222779, 260.336337731698, 258.520667047935, 259.178164538972, 
    257.408335627676, 256.484507173193, 260.507960894175, 256.945466922561, 
    258.127658176507, 257.779345626892, 259.115302610284, 258.575899148599, 
    256.796667112775, 256.977213365347, 257.874561137999, 258.196130927643, 
    258.418141343589, 258.11926150748, 257.660302542946, 257.142911997712, 
    257.942360636449, 258.423111931803, 258.566598228643, 258.972271511439, 
    258.832711221419, 257.342253533889, 256.842931400747, 257.497136177218, 
    257.468162568971, 257.549765243992, 258.337961164337, 259.363107878823, 
    259.11620354452, 258.557138106883, 258.448005415515, 258.651892278921, 
    258.212542530725, 258.820858073698, 258.766931176259, 258.738406023978, 
    257.366791898043, 260.131956113922, 258.517923896415, 260.243129554856,
  261.377934487574, 258.914803165012, 258.703135163185, 257.782754191957, 
    258.003699380187, 256.87275454357, 258.163228277612, 258.655037366269, 
    257.760849744915, 259.855099912575, 259.474060291713, 258.832687594411, 
    258.345063554264, 257.703430912598, 258.39746573636, 258.071009098256, 
    257.884926308239, 260.072104237778, 260.1329150929, 259.337043003719, 
    259.794230360145, 257.815627060482, 258.079483446809, 258.60250668531, 
    258.324543164068, 258.724723465417, 258.974149698173, 258.294230639635, 
    260.191711780957, 260.149381533373, 260.171453155531, 260.258775963737, 
    258.787700456998, 258.347498465676, 258.253498131387, 258.209638641317, 
    258.341236017313, 258.73185755592, 259.105254447919, 258.556580042528, 
    258.915528112201, 258.343664860683, 258.408155272815, 259.794926072815, 
    260.00503968562, 259.45374935452, 259.82710540888, 259.63450565798, 
    259.236954797681, 259.315474448138, 259.712318791177, 257.613137443621, 
    258.275758268885, 260.043298527966, 259.630610181015, 259.187244454115, 
    258.719216261254, 260.487641278102, 258.665604089361, 258.265468075,
  258.939523244978, 259.376108903558, 259.738226980307, 259.889827293536, 
    260.510703235406, 262.328644503903, 261.363573895406, 263.580526907558, 
    264.771994595136, 262.578827127531, 258.506804577013, 259.517808897814, 
    259.781791777667, 259.755865005546, 259.741061838361, 260.465307234864, 
    260.195233017462, 259.897564942122, 257.917962631255, 258.233234610652, 
    258.979035287051, 258.817734889088, 258.125357775684, 258.689359645281, 
    258.005339448425, 258.227827044219, 258.834043006592, 258.402967874259, 
    259.538873445706, 258.815817774604, 259.019226236092, 259.674750445621, 
    258.768664376403, 257.679572096228, 257.628160035197, 257.972591597306, 
    258.435942756206, 258.916562912623, 260.069760352569, 260.302367107983, 
    259.109518443902, 258.843456218941, 259.715124978389, 259.582645745579, 
    258.325528472052, 258.336293876057, 259.072230290128, 259.073597565972, 
    258.880370395414, 259.66161369846, 260.503930033371, 257.941495924219, 
    258.184247417791, 259.435629361068, 260.051091667385, 260.070471343153, 
    259.67192198553, 259.292032741929, 261.819862917607, 259.406009097077,
  254.369227075442, 257.050139623366, 258.576789226784, 257.86542347721, 
    257.478314734749, 259.58289420013, 259.456542915074, 258.080355452126, 
    259.837264246388, 261.724522412241, 260.434487136706, 258.765798443394, 
    257.515651683206, 258.009774283104, 259.355329572468, 259.209989858975, 
    258.767613113803, 258.035466958548, 257.672539190097, 258.387752375138, 
    257.528050917688, 257.096753169661, 256.693572460476, 257.563561068801, 
    257.565890185898, 257.724893726042, 258.794497804371, 259.963390914178, 
    259.922579462646, 257.032346952199, 256.051132205027, 256.844416656468, 
    257.812200937012, 258.356616814902, 257.801297664023, 257.464101624338, 
    256.991689960005, 257.440603522478, 258.438542719204, 258.634749303714, 
    259.396168842385, 259.410779794873, 258.777964673451, 259.115578196989, 
    258.426364289003, 258.108283194507, 258.452194238518, 258.227557087451, 
    258.547935537661, 259.136166070806, 259.116257706272, 259.033250750446, 
    259.304014765117, 259.320910645566, 259.74226349251, 259.146629080256, 
    258.823617324462, 258.567287182639, 259.822889473295, 258.282212543586,
  256.330287595541, 258.649849019068, 257.542857713171, 256.309057399216, 
    256.183711170698, 257.888567692765, 258.62215281774, 257.754655975738, 
    257.262826038663, 255.947017641659, 257.236624920135, 258.030030131305, 
    256.261574466033, 255.842089250716, 257.487017394701, 258.113082089163, 
    257.576428950189, 257.533729170808, 256.631364355223, 258.182228685153, 
    258.837137757626, 257.10809204809, 257.708420272314, 256.603558950383, 
    256.077614777047, 257.853029749096, 258.523283615449, 258.667446686972, 
    259.971995332234, 259.041745526838, 258.885369978615, 256.116203180746, 
    256.681279676145, 256.079890693787, 256.7656116917, 257.36681043064, 
    257.463561131612, 257.312413116995, 257.488165526772, 256.858302777064, 
    258.605823352632, 258.90544472459, 258.33288538102, 259.592920121531, 
    260.062391231584, 258.926650275966, 257.907119650509, 258.065909215729, 
    257.996682529946, 257.83036665967, 257.940728975823, 258.240950446505, 
    258.202751953186, 257.592186844395, 258.202279408094, 258.982127391782, 
    259.474578832749, 257.447050695274, 259.070903285468, 261.004288878023,
  258.446822925674, 260.664126157489, 257.664847218925, 256.521904641538, 
    256.257168350178, 256.576540331616, 256.414580503987, 256.045527270233, 
    256.831934008519, 256.001403828373, 256.130311602415, 257.786387154133, 
    257.899960746883, 257.01048052981, 255.689787403107, 256.870882978709, 
    258.630056370753, 258.624645335707, 256.102335353461, 257.048626881531, 
    259.318092704403, 258.665676318054, 256.921926227366, 257.51334221388, 
    257.451920337285, 256.994172449888, 258.553868816018, 256.884095541887, 
    258.523568919614, 257.66245474749, 256.912289823668, 257.159400786162, 
    256.877718296932, 258.111857377741, 256.876791024402, 256.938798829557, 
    257.86493503687, 257.722721173436, 256.21480047692, 255.147017469607, 
    255.266563028286, 257.289324798149, 258.79853440294, 258.890985351494, 
    258.510128041264, 259.008304356695, 257.655584931464, 256.362601434522, 
    259.02288855971, 257.355385481844, 256.931982581576, 260.14254732117, 
    258.524272273366, 257.749652094859, 258.29282908868, 257.754705980429, 
    258.101178913026, 255.157464986279, 257.721625575184, 259.288485875922,
  256.65369295618, 257.45830869106, 257.661145370474, 257.159905803173, 
    257.170116787611, 258.379805831647, 257.936979593821, 259.715861212002, 
    258.715053992391, 256.007333106519, 255.442547190702, 256.18420823091, 
    257.884399041953, 258.90526788119, 255.496171373098, 254.050234404582, 
    253.83524463255, 254.512761456661, 254.172853838121, 255.75628257106, 
    258.915132456029, 256.915683380871, 253.188518711911, 252.555419320961, 
    256.775413728014, 256.374129547795, 256.824695485269, 257.081697363162, 
    255.98451902552, 255.059141736269, 254.634148034785, 253.304697989211, 
    252.758752899543, 256.189052285632, 257.566500739963, 259.504059035142, 
    260.937034885558, 260.562656798036, 257.099523772028, 253.147622078627, 
    252.876977285282, 254.66714736816, 257.01391635132, 258.538403823975, 
    258.030135460464, 258.748496201153, 258.586065480679, 255.782091323343, 
    255.287484983426, 256.261064710975, 253.961641539937, 255.42213907188, 
    257.78211735777, 257.687232854818, 258.643891164255, 259.051520154483, 
    256.343041720166, 254.450842192113, 255.942801030922, 255.635703891088,
  252.414762724371, 253.942738158688, 252.5733518664, 251.77542413116, 
    252.823749460778, 255.418431110366, 256.854951262526, 257.57620233258, 
    256.731532297874, 250.779665613765, 250.212088575467, 252.338107521188, 
    255.147032786782, 257.12758541516, 256.897610087652, 252.925791810683, 
    249.805228144935, 250.623101174318, 250.51245811611, 250.757262807036, 
    253.922513122849, 253.151792594095, 250.122200964039, 249.252535756196, 
    251.574267894398, 251.695615503686, 252.461315402968, 252.936675054059, 
    252.424718199107, 251.700922797848, 251.742121662454, 250.029123479278, 
    247.472005650921, 250.262886188278, 253.2516444992, 256.15144753175, 
    259.177845968178, 258.304586447781, 254.199335176397, 249.872269463212, 
    247.745536935546, 250.29392507097, 252.685539475017, 254.096044899518, 
    254.7127105299, 255.211882080382, 254.597873262058, 250.8593584202, 
    248.662111071554, 249.902888028865, 249.358436806961, 250.167548606407, 
    251.65859418791, 253.17851749219, 253.923298938856, 253.454553405891, 
    252.577756331126, 249.710883045557, 251.036871191438, 252.215298483371,
  247.690382673578, 248.114792406901, 247.883043444228, 247.897036562113, 
    248.030874377362, 250.077737469982, 250.566032386091, 251.171242921985, 
    250.385873951906, 246.330272666242, 244.609972223075, 248.221810212829, 
    251.026889588442, 253.278069316928, 252.429030535244, 249.075059805189, 
    246.431442743814, 246.812460388178, 247.095696443181, 246.959476731882, 
    248.383317797203, 247.845570375041, 247.695208612787, 247.042113792597, 
    248.514040432792, 247.767757760754, 249.304233438059, 249.203394933608, 
    248.730939975113, 248.827857439724, 247.35082951781, 245.484657338024, 
    244.300818792308, 244.991706917827, 247.740581274539, 250.148698378578, 
    253.418155219479, 252.490660350848, 247.429637768995, 245.488869379503, 
    244.489398279639, 245.622577016596, 249.058126258457, 250.182700629206, 
    249.768526143613, 249.905833000648, 247.725507164276, 244.886895077664, 
    243.338153973117, 243.954886412844, 243.884932799211, 244.286550301299, 
    246.238947346628, 247.444400607065, 249.678428318962, 249.952152756525, 
    247.7023966093, 246.620881658114, 244.599207338534, 246.297254369854,
  242.348264400088, 239.719000292869, 245.070180693007, 246.849315818661, 
    247.04828129911, 247.551795448903, 249.330975186176, 248.944588660685, 
    246.566881239518, 244.878786267584, 243.213707877476, 244.809762588507, 
    247.097823557662, 248.502228684138, 247.825338027196, 245.614838492793, 
    242.605539733734, 242.413764686869, 243.850751818517, 244.878178639973, 
    245.911358793242, 244.884012178269, 243.935952825797, 244.540007014162, 
    243.680894347494, 245.751784442141, 248.980420598658, 248.371769733392, 
    247.480449838969, 244.670838497949, 242.623754246403, 242.552319788441, 
    242.39290077294, 242.954451573609, 245.774860467841, 248.367698730107, 
    248.77304189245, 247.039995601959, 244.062134919968, 242.968090811459, 
    243.571213261829, 245.163468508075, 247.332776767902, 247.453615546633, 
    248.840688250005, 247.906445831929, 244.405803899383, 241.907759167997, 
    240.905452435624, 242.027420343823, 242.412616370436, 242.294279751769, 
    243.487425836191, 243.065723502543, 243.665168116766, 246.785665691821, 
    247.818498906696, 245.07087829043, 240.817670762365, 242.802884692342,
  239.431168475653, 245.08988993562, 246.057575986909, 244.519053943794, 
    245.408982887174, 245.512636667134, 244.239864618179, 238.931259122165, 
    237.243299031601, 241.261495757534, 242.596237435903, 243.350653467629, 
    244.183591526358, 243.257242293332, 241.633377411948, 239.329518340409, 
    238.530881657229, 238.506071377531, 240.308212989653, 242.554743225262, 
    241.795335796879, 237.978152975434, 240.776695691425, 245.599691688189, 
    245.530747862322, 246.171668010663, 244.250690816995, 243.364358674496, 
    242.41217792247, 240.220673951437, 240.691381344824, 242.096592539452, 
    241.765818654357, 242.071001363584, 242.838209031088, 241.978308747233, 
    239.097284856874, 238.181861251367, 238.014829318608, 240.223105014381, 
    244.752238560212, 246.345647278215, 246.744507352966, 247.239682937319, 
    244.814416196158, 241.799094236008, 238.87284500222, 238.624475493048, 
    243.33873283831, 246.340450000654, 241.928451615458, 244.07202276558, 
    244.635098837411, 244.687997721041, 245.649777592609, 247.069427690624, 
    246.117732643079, 241.11005345789, 238.623329725393, 237.315352867879,
  237.308214832458, 241.565981565977, 241.971154570983, 239.771848898972, 
    239.031525678883, 239.353565493267, 239.670534870886, 239.498621966175, 
    238.999914683945, 240.447084917138, 241.018274894297, 241.323420015363, 
    240.711935434694, 239.249207746911, 237.90997259891, 236.673210951524, 
    236.339718371543, 235.346771315985, 235.825546879117, 239.104218845297, 
    240.317032042148, 241.627987751077, 243.750468682686, 243.368663279896, 
    241.493908791021, 240.288313228573, 239.939777850755, 239.762239007094, 
    238.170199830361, 236.737500980544, 236.413000979374, 238.171960744702, 
    240.972917326409, 241.582821240183, 239.920121988386, 237.714277732615, 
    236.848895262733, 236.027597333106, 236.90953704692, 233.923463254413, 
    236.632417700152, 242.05705403285, 242.628219552047, 240.656319817774, 
    237.669722961847, 236.02642883441, 237.981208011308, 243.336840791175, 
    246.600631950934, 242.558736220641, 238.871186219199, 239.778353567576, 
    239.566862511669, 239.923810752963, 239.188737195772, 238.581317459302, 
    238.254494196847, 238.172162682033, 237.751103791319, 238.576231083067,
  237.624916778552, 240.069841347941, 240.776003719535, 239.423452280075, 
    238.277332001205, 238.106732678053, 237.868186513347, 237.246649951699, 
    236.609732440013, 237.93995979369, 239.860613676754, 240.613723021084, 
    239.430200710453, 237.669699569523, 236.882067761818, 236.183174161405, 
    235.321201277596, 235.224043875868, 235.738032266551, 237.381094504904, 
    238.589656831759, 240.235702078078, 240.74957581073, 239.415348832025, 
    238.793190498507, 238.756764067457, 238.214594025784, 237.541118692551, 
    237.021435877381, 236.359596312321, 235.470008546953, 235.123505292986, 
    236.212335407575, 236.53863746394, 236.401299889042, 236.350811352111, 
    234.578271715727, 233.337555622603, 238.738917674707, 241.436516213327, 
    241.835177808321, 244.903231369967, 244.175578412242, 242.554471583068, 
    242.593695891443, 241.483311672714, 240.088707627174, 238.752451361452, 
    238.80972224977, 239.5014983642, 239.45374369195, 236.88542625241, 
    235.648181527887, 233.945119593311, 233.357371905095, 233.772811171305, 
    234.585956734245, 235.389892163993, 234.68030937094, 236.184993857023,
  232.55446767609, 233.763523866352, 234.655478196065, 235.026568332012, 
    234.835912480865, 234.18952983097, 233.458043244314, 232.531485444854, 
    231.78156916518, 231.948776370369, 232.846292685466, 234.100128282534, 
    235.091068897858, 235.152981419386, 234.995472436697, 235.364352381977, 
    237.871212562777, 240.040239116725, 239.367500992871, 239.324871210201, 
    239.022360412406, 239.114323255233, 238.981173460595, 238.838026558687, 
    238.909887449997, 238.826799939495, 238.127231691229, 236.987374957964, 
    236.108400647939, 235.372825806101, 234.43327995799, 233.702450857303, 
    233.955525680353, 234.692184386717, 234.907293553045, 234.574055626697, 
    234.464409977798, 233.700747868158, 233.012285602658, 235.976597249046, 
    238.671319327181, 241.762522657088, 243.195061526712, 243.650020802532, 
    243.978937127286, 243.13596100845, 242.337467494843, 240.328595999325, 
    238.210886837801, 236.879290927694, 235.429162572206, 234.499733857286, 
    234.683300182103, 234.049972495762, 232.926621567288, 232.083328357767, 
    231.05350851497, 230.774627770635, 230.56381323752, 231.430291684078,
  228.812065209852, 229.156393366438, 229.612789212557, 229.819273909662, 
    229.800687591249, 229.731768804017, 228.949560381829, 227.777607235034, 
    227.325430103502, 227.612898289478, 228.275028932025, 228.943674362093, 
    229.421581947531, 229.91535009213, 229.923846668392, 230.668489084122, 
    230.928667062987, 232.015761097621, 233.240122811126, 234.342464575092, 
    235.26390829051, 236.130110683549, 236.857780744128, 237.409139010432, 
    237.55701618731, 237.53668568171, 237.107312834128, 236.432481632822, 
    235.987974282361, 234.687712064268, 232.579898443891, 230.968388394781, 
    230.538542880106, 231.008284052464, 231.584969519183, 231.812962357023, 
    232.35056920613, 233.645370437742, 233.558987963111, 233.016729768438, 
    233.582181595179, 234.50152348388, 235.127586341026, 235.381053319007, 
    235.03659026517, 234.555228775168, 233.865636545271, 232.562040872528, 
    231.187303705259, 230.281053261835, 230.133808952833, 230.724350182845, 
    231.759293470102, 232.386189761336, 232.150423707112, 231.260899784474, 
    230.015591801589, 228.895556925129, 228.672188479971, 228.707847749952,
  227.042475865825, 226.941544084268, 226.746294496255, 226.533520791785, 
    226.217104016191, 225.764204350149, 225.414661234914, 225.300072986787, 
    225.217417293937, 225.277747777117, 225.599521900712, 226.078751703027, 
    226.595077250867, 227.050938175207, 227.487848139014, 228.086814960193, 
    228.373641385386, 228.814075638082, 229.204215988511, 229.724828229332, 
    230.371913660003, 230.998421345828, 231.37268666382, 231.772091606528, 
    231.961834438145, 231.858926714773, 231.664712071431, 231.0594365775, 
    229.956396203356, 229.134657681809, 228.636708747406, 228.237619514149, 
    227.850822390778, 227.640002767919, 227.674641963619, 227.814863272461, 
    227.95354875154, 227.760994097156, 227.223333279073, 226.738702860394, 
    226.397565405468, 226.324629771496, 226.5765619483, 226.933876631488, 
    227.216515270069, 227.367387568138, 227.558093092417, 227.754411967973, 
    228.0269238608, 228.372498321059, 228.730955786514, 228.999170223131, 
    229.098938839513, 229.301457526695, 229.431031760418, 229.224749846426, 
    229.224371221893, 228.712571870995, 227.454819821579, 227.024483649528,
  225.180892674757, 225.378493398316, 225.742964838867, 226.099143743913, 
    226.225664729966, 226.24407068579, 226.233660575673, 226.30358459739, 
    226.498912307728, 226.834847953246, 227.15230865634, 227.289872906274, 
    227.238443647938, 227.088434117121, 226.941600105866, 226.66548984861, 
    226.245093756677, 225.771413651587, 225.378035467776, 224.969350121803, 
    224.603905834589, 224.287581016945, 224.095987012405, 223.983459280409, 
    223.977751558362, 223.9084851157, 223.822196017415, 223.732775906535, 
    223.509640288821, 223.068083578357, 222.961468439826, 223.624989997454, 
    224.834699998952, 226.00639503306, 226.736613895027, 226.964136761895, 
    226.810311338551, 226.521855499616, 226.295055697061, 226.069480504047, 
    225.893732397905, 225.823155985115, 225.703143952096, 225.475025227814, 
    225.197911077086, 224.945752565528, 224.680457239482, 224.379404496235, 
    224.079879370584, 223.934914647532, 223.898708516988, 223.953859448643, 
    224.002048270189, 223.850588150608, 223.474575055727, 223.040505291444, 
    222.7493055571, 222.802636193482, 223.605310163459, 224.659411298948,
  248.022636120453, 248.061395928634, 248.034465822615, 247.872256099813, 
    247.629514290013, 247.365118439515, 247.219466203548, 247.038754265053, 
    246.845904760222, 246.523837360817, 246.167471307436, 245.867291647122, 
    245.649273443688, 245.435391960069, 245.379297279302, 245.326210798919, 
    245.420603341761, 245.66974610261, 245.594415930976, 245.700605407125, 
    246.286970674241, 247.124833275057, 247.700051327407, 247.790971322758, 
    247.421877523128, 246.865750406447, 246.581303085021, 246.723271515931, 
    246.887259708954, 246.90927488062, 246.769428455726, 246.432780959359, 
    246.377990781002, 246.562659708815, 246.770639135306, 246.988957064396, 
    247.224716898795, 247.362769503819, 247.429838249104, 247.481896167579, 
    247.538384649649, 247.61838546789, 247.722504457132, 247.789085460941, 
    247.784771622609, 247.70088476811, 247.655522184671, 247.647883795902, 
    247.59904794696, 247.547056493055, 247.512470644467, 247.536011879309, 
    247.57053126605, 247.622476844029, 247.69169836225, 247.73826298228, 
    247.813180467361, 247.902695721664, 247.974026154108, 248.010071858151,
  252.782049783117, 253.068258247748, 253.352893895275, 253.201824057702, 
    252.417812184271, 251.327655599814, 250.374448794387, 249.676970262179, 
    249.029187683006, 248.278261982072, 247.337008121471, 246.712964973463, 
    246.452253804385, 246.471138459464, 246.784668209489, 247.138265002614, 
    247.37641259807, 248.025255973692, 248.635429694007, 248.621684606761, 
    248.120764439045, 247.905016582109, 248.139411583941, 248.197746559901, 
    247.740983788996, 246.866467370134, 246.156668861373, 245.696528877811, 
    245.325691321145, 245.321741412563, 245.721609580431, 246.334631571658, 
    247.21026202775, 248.095680362229, 248.592781523389, 248.99375789192, 
    249.456175591363, 250.005194855507, 250.309314332022, 250.702586886421, 
    251.026820127358, 251.07848688444, 250.832056416038, 250.687455184236, 
    250.620075412425, 250.273416157348, 249.971904902172, 250.07765391454, 
    250.277142981522, 250.380880393709, 250.508551044126, 250.664858292805, 
    250.879438860236, 251.082830024944, 251.364425267133, 251.614198090752, 
    251.784617851932, 252.096888295433, 252.403525712851, 252.621481251138,
  254.473296465754, 253.950862979634, 253.664136129095, 253.118634871854, 
    252.613218943642, 251.926732309214, 251.200950873111, 249.783300107852, 
    249.043921916807, 249.993371551704, 251.323829575629, 252.397537816053, 
    252.529905459275, 252.369681102502, 252.290516670684, 252.379404627582, 
    252.672723146393, 252.466025838776, 251.707885855634, 251.728863690579, 
    251.326508545953, 251.685246241388, 251.263263338364, 250.442185679468, 
    249.255453633629, 247.739076161874, 246.778266892607, 246.912991828895, 
    247.707642840079, 248.581905134694, 248.998886602279, 248.846928699532, 
    248.806336254644, 248.955179944903, 248.769570899153, 248.54948962468, 
    248.667318503323, 249.503935282073, 250.611884715274, 252.147035212295, 
    253.679640862437, 254.592130345354, 254.321730449071, 253.399718595311, 
    253.05352137824, 253.222773284338, 252.977844274257, 252.0008839407, 
    251.113302188446, 250.604571447514, 250.282052961363, 250.009486380807, 
    249.800283190928, 249.470313472261, 249.449824604718, 250.201067670829, 
    251.063806869505, 252.276811881817, 253.578178106528, 254.473463458807,
  256.17013078491, 254.801577496124, 253.332886643929, 253.370963770719, 
    253.826579054251, 251.822470678182, 250.142340035625, 251.958887592365, 
    255.00457884454, 257.560704477207, 259.619308903293, 260.29306210058, 
    259.894468592905, 259.426066600999, 258.270751521268, 256.022271935965, 
    254.644535452752, 253.461994096643, 257.2369712033, 259.493891218709, 
    260.040857035374, 260.91351687333, 261.228117698332, 259.673509029179, 
    257.186791245243, 255.594854604588, 253.51409227078, 251.90936078138, 
    252.253625945121, 253.176879256736, 252.691608277882, 250.404942401475, 
    249.108399851478, 248.6314912901, 248.278098885543, 248.44005005491, 
    247.70902015953, 247.934861552231, 250.923576217492, 255.297920482795, 
    257.684370308754, 258.410403213647, 257.96623823697, 256.098582995792, 
    253.799040751374, 252.171636910942, 251.209910906729, 251.28184568264, 
    252.339664922787, 254.566543756408, 256.31215023968, 257.502570069919, 
    258.004494212297, 257.902959347009, 256.813880106698, 256.32855917769, 
    255.56827661753, 254.966105426114, 255.603323628868, 256.558353934994,
  261.303983290325, 259.731338171271, 258.529569370928, 257.045356063782, 
    254.712957537784, 252.587804427244, 251.871885171221, 255.508721333714, 
    260.582857937467, 263.148768868696, 263.650886203027, 262.630556359557, 
    262.281200028908, 261.339038214815, 259.68246758599, 257.624969767451, 
    256.651975819417, 258.441882623387, 261.859120514587, 263.248057574733, 
    264.575377357956, 264.550123764996, 264.059455332632, 263.865781807542, 
    263.304082295963, 261.066710048505, 257.808762309944, 258.021033581859, 
    256.248680318218, 252.47468655598, 249.960283755257, 250.322860118279, 
    250.632733494092, 250.638649729262, 250.933671461932, 250.374377190618, 
    248.969824595417, 252.475985928676, 258.273846760174, 261.391912331661, 
    261.183167311947, 259.724676585217, 258.798234297892, 257.080667999283, 
    254.661785694677, 253.732450253709, 254.39426861914, 255.295924959051, 
    256.554879418984, 258.502929629868, 260.415531394903, 262.963290358809, 
    262.398272755131, 263.684874176138, 264.941554388557, 261.881766516358, 
    258.653568350688, 258.718085080781, 260.116123831864, 261.760347670217,
  261.489818375909, 259.563503135838, 257.54653861246, 256.336668335566, 
    255.712878180052, 254.498302882783, 254.851653020811, 257.606810231287, 
    261.643259855508, 264.332462185176, 264.216832871445, 264.592887619034, 
    264.527913211762, 264.380494386729, 262.077398029032, 256.243356871836, 
    258.30767000895, 260.291656757578, 261.61870360236, 263.745667881178, 
    264.7586835989, 264.846983716784, 263.84475834167, 264.001554760778, 
    264.040433307966, 263.926209815661, 262.466662246792, 258.609636625588, 
    252.646287331565, 252.415558754511, 256.131317269864, 258.270610971471, 
    260.606411996182, 260.617609456994, 259.212787015757, 257.487907676655, 
    256.559541600344, 257.8600017534, 259.876802820617, 260.812249417815, 
    260.917580759398, 259.536703280264, 257.605070922776, 255.904086985477, 
    254.945469063401, 255.434545537808, 256.61518806643, 257.617204985925, 
    258.057645793353, 259.17346199979, 261.638877415202, 263.194335552754, 
    262.724132304757, 262.881122542273, 261.727104215615, 261.330057846259, 
    261.624428557447, 263.286507736135, 263.597466667023, 262.389568452127,
  263.045691013656, 261.262585380437, 260.033628198551, 258.093166360641, 
    257.637190530181, 257.687653579114, 258.473087925831, 259.573480232844, 
    262.430804008136, 265.348253116707, 265.670825801674, 264.457001513268, 
    262.657491441941, 264.26808207534, 264.163188865826, 260.092687726286, 
    259.204902048058, 261.498567657826, 263.520626918097, 265.887316446739, 
    265.949315275428, 266.440226641729, 263.360964697708, 262.11671251683, 
    261.120277780207, 260.404524049593, 258.774363879032, 255.106689703287, 
    253.703977389687, 258.916579586567, 262.011954449461, 263.774857191723, 
    265.179933134609, 263.47460310981, 259.886319281956, 258.039365071936, 
    257.038783636617, 258.142919870263, 261.465758122423, 262.759391060481, 
    262.801790399724, 262.091328696799, 260.699479365249, 259.559097069591, 
    259.467097381475, 261.171927251777, 262.631051251452, 263.459212949015, 
    263.452449868234, 263.202101620125, 262.776879987013, 263.474726264357, 
    263.625936160851, 263.306281077231, 262.123286589641, 258.515827610854, 
    260.518421521673, 262.182253425325, 261.042682198557, 261.871755253491,
  265.343489430133, 268.36999891912, 265.87509644533, 263.511591954917, 
    261.005245162141, 261.808543996201, 262.915230321859, 262.437262844192, 
    263.197700118155, 262.955910828348, 263.787940619466, 268.13335184791, 
    263.531038751865, 262.634164114114, 262.260877123712, 264.641708155836, 
    263.623159022445, 260.196162510645, 262.979464908363, 266.722329427262, 
    266.947026531486, 268.739238466927, 267.439949324625, 264.546897399262, 
    260.820258094928, 259.099545024458, 258.294729055683, 258.66256764882, 
    259.606072922257, 261.308401206264, 264.066917643437, 265.115903947118, 
    264.463921541791, 264.987689358734, 263.370931977175, 263.218535243903, 
    262.438705265381, 261.812984855485, 262.1711256021, 263.291212529036, 
    265.349677334046, 266.105602188833, 264.947764580928, 264.286209540918, 
    264.428479048575, 265.290342501623, 266.01590500175, 266.598679541244, 
    266.825054980574, 266.72634104192, 266.821192363476, 265.042797584866, 
    265.753690053544, 266.359471480304, 264.042745553059, 263.449307617737, 
    261.473623779204, 258.362533666604, 258.443521446454, 261.527296255376,
  265.812461090875, 268.166281041727, 268.600179614342, 265.952309065276, 
    264.20302851242, 266.29147860514, 267.469514599369, 266.583974551452, 
    267.174570897392, 267.766076213291, 263.378193141281, 267.072736087829, 
    267.486287696715, 264.43431927096, 265.895880629671, 265.800620507567, 
    268.546904767997, 266.072718716509, 262.540102826558, 261.277847787745, 
    262.869363577671, 265.339865472332, 269.124553717706, 270.165109794191, 
    267.158668987574, 264.182414364228, 263.647848439763, 264.976944758634, 
    268.56498458074, 269.57574677299, 270.066337302257, 267.220409411002, 
    267.168033006308, 268.769867565502, 268.741845243601, 269.260584345684, 
    269.349634453328, 268.79011405319, 268.287320263158, 266.96167485509, 
    266.589511548971, 267.344805681992, 268.334027877151, 268.209997110594, 
    267.053439944563, 265.799067987957, 265.724829253065, 266.318518902349, 
    269.089472942485, 268.824673761746, 269.501437705117, 269.44527692195, 
    268.76763534758, 271.399482281714, 273.665722261086, 270.930885627428, 
    268.107765853791, 264.498867067684, 263.840506777229, 264.368711786408,
  272.71530525097, 273.698209614364, 272.25775734165, 271.136473517954, 
    267.651120630936, 267.970750825556, 270.510905498095, 270.993177533889, 
    270.808560758278, 271.647333774053, 270.18487767906, 271.906742741427, 
    271.587637485685, 268.008479559817, 270.692784732214, 272.914933625763, 
    271.295088416076, 268.419696362696, 265.814685477612, 265.893384317135, 
    265.433667182496, 267.110348248797, 270.656141411066, 270.846801598713, 
    270.625105269158, 267.992135980101, 265.400003068666, 268.187802264061, 
    275.408322498268, 278.088698568064, 275.512198932852, 271.004643243616, 
    269.775054726833, 269.677070331264, 266.134869214209, 268.420260029165, 
    274.038697147984, 273.695423644836, 270.633632360167, 269.07255571478, 
    268.465005185507, 270.387030835614, 271.915627100407, 272.487022795965, 
    269.92813478885, 268.359094507407, 269.890303786826, 267.872963144517, 
    269.611412365497, 272.432854830738, 270.826089910733, 271.015506408981, 
    270.977773819645, 273.63021076152, 275.977953993264, 276.349380270655, 
    273.394407853433, 270.28928815658, 267.367305167618, 268.239386611844,
  277.387140381198, 278.423583641046, 279.617679122611, 277.230704150376, 
    273.454079264061, 274.896091920633, 276.630826829857, 276.443829942111, 
    278.573519753709, 277.171331846639, 274.471802694311, 278.029713846081, 
    278.668995420989, 275.777539124332, 278.891232745843, 279.786389480187, 
    274.235751548673, 275.250492031072, 273.556023923033, 271.547980200597, 
    271.123386194123, 275.511150712629, 280.55109662275, 276.958528191003, 
    273.317350813461, 267.504629145265, 267.931847953286, 273.674988073782, 
    278.233719123819, 280.551283558716, 280.555876751799, 279.170482807, 
    277.378454426391, 274.045467474022, 273.806590405314, 276.624476739935, 
    279.145206017801, 279.70351391129, 276.844026478372, 272.015366294084, 
    272.018442494776, 275.46975186881, 276.713475061931, 277.905877173141, 
    276.390560693443, 273.557740063316, 271.718248118609, 272.362433671925, 
    274.037643084291, 277.515491385754, 278.201747983854, 275.858558131961, 
    273.330560530869, 274.230250457712, 278.488867440285, 280.803075828871, 
    279.032648733512, 276.411648258437, 271.542720610917, 273.165293716101,
  282.627974086121, 283.80221567769, 284.8706992122, 281.811211068902, 
    280.657036271262, 279.296330059666, 279.739313171879, 280.9070766858, 
    277.954758649397, 278.475361211602, 282.459708037164, 283.166491305907, 
    282.42027889979, 283.65995720353, 284.279217003342, 281.114006246203, 
    279.453547603893, 278.269054969435, 277.581347879462, 280.544766734917, 
    283.016522679855, 285.064263300301, 285.077982083421, 279.471734690153, 
    276.758886658744, 274.671905923328, 277.868888456451, 283.045290750929, 
    286.823814935334, 285.496941617347, 284.569995216732, 283.136449275724, 
    280.248144546805, 279.4234655461, 282.977307760737, 285.623540156543, 
    283.937134929187, 285.158609843595, 282.896698528112, 278.269040475559, 
    278.909819584217, 281.913760108118, 282.653406579241, 283.680174776427, 
    282.114908251961, 279.696765955707, 280.04599883548, 283.726250367471, 
    283.279389546788, 282.184766407439, 283.680488534308, 281.468856727159, 
    280.098578785663, 282.480675046496, 284.636043412084, 287.20634742329, 
    285.096042351404, 279.746604979345, 275.703592667652, 280.082410221823,
  286.654972919044, 286.919523541177, 284.815885348124, 284.198637212934, 
    282.96782207861, 282.404600806276, 282.247701524527, 284.347188051992, 
    286.084426054885, 286.586206609845, 285.840252732564, 285.290106282801, 
    284.715479891485, 284.759337642041, 284.570721071448, 285.425354739653, 
    283.692667804536, 281.374509686032, 283.257194810554, 285.22597702417, 
    287.83329152346, 286.744093217975, 287.992878148489, 286.648907852405, 
    282.936255764362, 284.349829569715, 286.115698840139, 284.949168187531, 
    286.175197828478, 288.010020720876, 286.746258161299, 284.444240420462, 
    284.184967289445, 285.734780240204, 284.804438498763, 285.498523766378, 
    286.019426943866, 285.369319907969, 283.755009763924, 281.813786525494, 
    281.793979243723, 285.575543710797, 286.89400544754, 284.69829547092, 
    283.060582537532, 284.090250038192, 285.204143306431, 284.396722723703, 
    285.240028712496, 286.973604173964, 286.583559885427, 284.698371683522, 
    284.423678118031, 285.845404084537, 285.613852020309, 285.094158088875, 
    284.703732898112, 282.018600264136, 283.063445304934, 285.961312452507,
  282.796361638958, 285.350904312992, 284.313412549463, 283.92360482614, 
    285.184461182453, 286.9049965215, 285.481342310804, 284.776822680874, 
    287.110523952991, 287.089099211902, 284.229696196714, 283.93333193204, 
    286.458062222931, 287.206646962995, 286.50349238025, 285.631775054468, 
    283.558267595411, 286.081765533233, 285.740919065346, 283.47995360208, 
    283.709651509238, 286.27382017931, 287.762696942758, 286.912204545782, 
    287.293607862667, 285.170577334581, 282.613386452492, 284.90733247384, 
    285.294008224014, 286.035239859303, 285.358837832897, 284.580901232579, 
    283.68556809324, 283.705587453941, 285.42468158147, 285.560455547503, 
    284.710357036062, 284.276914814998, 284.251128150009, 285.474340168861, 
    285.04519308036, 284.997250353281, 284.512061301292, 284.104132460534, 
    285.001356631631, 284.39505236296, 284.069570438271, 284.419888984328, 
    285.559442866186, 285.232979042661, 285.415247917993, 287.040866771517, 
    285.446244904368, 283.850028448011, 285.40132926606, 285.894750464229, 
    285.713742840026, 284.097585418176, 285.051098615384, 284.65279516075,
  282.511302204743, 284.274906349962, 284.834625709596, 285.949201060517, 
    286.791993453499, 285.891674744395, 283.461054044065, 284.899139465501, 
    282.335706877091, 282.206309530007, 283.106444431503, 284.351998497086, 
    285.376016547723, 285.891410803778, 285.579431624902, 285.941227306173, 
    285.125290545986, 283.325346031742, 282.953988431598, 282.109587765203, 
    283.333195069272, 285.532843035117, 285.952324644297, 284.402708415898, 
    283.487968585129, 283.35880898448, 283.699580864042, 283.889593880974, 
    283.106771100929, 283.5186538426, 283.20620377927, 282.25570982144, 
    282.844249604176, 283.073346827266, 283.720039224509, 284.565571256127, 
    284.508140399875, 284.108614207339, 283.661729674564, 284.381206274059, 
    283.99415240135, 283.999166866538, 283.476774520143, 283.162217683844, 
    283.250289689331, 283.015198688968, 282.840455919437, 283.469910620933, 
    284.35434584782, 284.368122336973, 283.213339468407, 285.330447416101, 
    284.645854083771, 282.874032365901, 283.638968952983, 284.143939168982, 
    284.167479887137, 283.386576728339, 284.844427076359, 284.542333203837,
  283.442273171732, 283.031729083276, 282.923308623087, 283.395350069567, 
    282.317104997256, 281.283481078608, 283.549833706691, 281.367899826799, 
    281.017787304932, 281.51883138319, 283.1373929984, 283.192135305813, 
    283.110726136242, 283.199903548389, 283.068387120795, 282.068174354947, 
    282.401364817194, 283.322706353945, 283.698766728349, 284.356763777177, 
    283.10623669317, 283.776163320222, 284.040262077804, 283.11717204785, 
    284.12172262161, 283.221247368174, 284.352999508244, 285.05294601332, 
    284.137342362182, 284.997442778203, 285.187739719894, 284.115293174713, 
    283.139623655321, 284.098168105427, 284.89340629013, 283.97399119765, 
    283.478615806303, 283.491047880402, 282.3030055212, 282.593849680009, 
    283.820931566861, 283.708777002095, 283.064197804241, 283.446422546063, 
    285.525229115508, 284.787985901666, 283.843264053538, 283.633590247785, 
    283.627212911475, 283.650848497697, 283.398592125329, 284.445644793153, 
    284.362808250637, 283.098786081883, 283.22681650526, 283.339330682296, 
    284.107778051324, 284.815128571165, 283.843026032398, 284.836270503587,
  282.242777509953, 287.01206441674, 284.101776569751, 284.016999361061, 
    283.859494969633, 283.024044146744, 284.040152582174, 283.806155719057, 
    283.47426916478, 282.883334495542, 282.637931578598, 284.501713024292, 
    284.915487162084, 284.274023239075, 283.524163683673, 283.538693994022, 
    283.836518505893, 284.293231746069, 283.857201293524, 284.70253647757, 
    284.892387715387, 285.919438362081, 284.778516456315, 284.063258485901, 
    285.000866789468, 283.851533377522, 284.456249132916, 284.715458305814, 
    285.835191586322, 287.502307317982, 287.290851770754, 289.029430397296, 
    286.054318622016, 284.538588485736, 285.46337573888, 285.232449207518, 
    284.400441556284, 284.401876104423, 283.619061807714, 283.40157254991, 
    283.593759318454, 284.741528344256, 284.650004040402, 284.378996663835, 
    286.246084410544, 286.424042265394, 285.587946404358, 285.223188655275, 
    285.334605055542, 284.74167782934, 284.571850919001, 283.885635446217, 
    284.15112398734, 284.257405766641, 284.528441241311, 285.013104851945, 
    284.816685233335, 284.30334031001, 283.822935294825, 285.913081987638,
  286.627570331705, 290.185641048347, 285.195104853303, 285.937659933861, 
    284.507547042163, 283.393035007873, 284.833659962194, 285.279178058171, 
    285.009931960151, 285.112574703537, 283.459457666128, 284.665656577741, 
    285.301497646668, 284.124772369797, 283.557694064834, 284.305374708625, 
    284.167004576877, 283.918542347599, 283.541645837713, 283.085936612349, 
    284.674846888946, 286.329168609669, 283.965730829237, 282.556626929523, 
    284.225384432043, 284.166246765746, 285.73283164845, 285.311983761221, 
    284.120969683655, 286.015444620374, 286.2795239419, 285.399585378983, 
    286.471545226116, 285.06927364388, 285.239350969148, 284.295969293717, 
    284.224472218965, 284.023271458626, 282.374853613602, 281.823814230671, 
    281.496487764903, 283.400223513929, 284.408485505596, 283.889588702048, 
    285.924390258938, 285.937602402105, 284.823512522924, 284.326114118671, 
    284.798760036083, 285.545748564638, 284.911218860541, 283.19904154883, 
    284.007442203764, 284.63837118134, 283.594211274256, 283.7394903176, 
    284.759085036135, 285.977334865288, 283.757905441427, 284.882344331052,
  282.170822748535, 284.885941936634, 286.949296111491, 287.298011200861, 
    287.093358639409, 285.204400254918, 286.592848672172, 286.72445369186, 
    283.756662155585, 279.507166549915, 279.998765095939, 281.445415288849, 
    283.242278992856, 283.574824174873, 282.017803487997, 280.985923609105, 
    281.92536572882, 283.390560396774, 282.772806845747, 280.701128061532, 
    279.957320370411, 283.360863072836, 283.993652755959, 281.148540035385, 
    281.030029130399, 281.234316022652, 280.805792782209, 282.251838322448, 
    280.609292495427, 279.736302609482, 279.215526810633, 278.851236278606, 
    278.804429680892, 282.437190325368, 288.077967407855, 285.762313865612, 
    283.538858316908, 283.451738381707, 280.983397298697, 277.754942353298, 
    276.830295711526, 280.538657457082, 283.638443420868, 283.750138722074, 
    283.457110457277, 282.652631960185, 280.943361414812, 278.733385742888, 
    280.61919716674, 283.706384586448, 283.289926927537, 283.2637319728, 
    285.023301725209, 285.251031424175, 284.364906920533, 284.325942432708, 
    281.631741449976, 279.134827209512, 278.274921563429, 281.767061971614,
  277.56709353835, 277.42128077175, 277.490264859269, 274.813203828064, 
    280.08179699875, 283.133613089726, 282.437546760395, 280.848411712034, 
    278.740737313042, 273.716823296227, 270.97558531161, 277.128502387939, 
    280.981172127747, 281.417144493095, 281.287513703584, 278.963192263349, 
    276.034211513518, 276.569954292559, 279.861684285835, 278.858643636644, 
    279.738884817628, 280.474033184033, 278.625524459823, 277.04124544627, 
    277.792652841949, 281.333716669998, 279.112232098524, 277.876838546167, 
    277.684918074955, 276.386773232047, 273.750363733472, 272.430659274315, 
    270.709711435907, 272.518677365812, 281.206470482183, 283.560636034078, 
    284.217129216153, 284.868048439566, 279.728648932421, 273.44478259102, 
    270.081302535071, 272.703014727636, 277.749743869265, 280.220728197659, 
    280.532429529689, 279.362927726285, 278.378846282974, 274.945085925134, 
    271.553781426368, 274.280362617763, 277.737319475149, 277.681116388824, 
    279.275317418924, 282.242132834369, 282.234470553225, 282.126526551505, 
    276.770314870233, 274.199473021637, 271.04828193435, 275.004339234929,
  271.481484826114, 270.039389888753, 270.26337857845, 268.220708728709, 
    271.171756481545, 275.097911289431, 276.99284010281, 278.320464029523, 
    273.571789738989, 268.370568328386, 262.654972413438, 267.898536772374, 
    276.349079012237, 276.373683124107, 277.045393613211, 274.425332151388, 
    270.595529635559, 268.868142557129, 270.306763913236, 272.851331662843, 
    272.498323424051, 274.640835553385, 274.08768095877, 270.430868047492, 
    270.702345096731, 274.10595671427, 273.080617485029, 273.416549040691, 
    275.152577163702, 273.434493668235, 270.876114494213, 270.031820432404, 
    267.626092855177, 263.681097054027, 268.913632799449, 275.67491325489, 
    278.532825440773, 277.134928712246, 271.934434808763, 267.673169837697, 
    265.716495091866, 266.169955681778, 268.277815683228, 273.393043963611, 
    275.657283495165, 274.679111551318, 272.765405720401, 270.590896585257, 
    267.550652467409, 267.154129696281, 266.939731349092, 267.903485097318, 
    271.233533342144, 274.866986237318, 275.046440233962, 277.186405509846, 
    272.263405414712, 268.558262328878, 271.494373710081, 273.430505615641,
  264.756703748984, 264.157358396412, 265.996800160644, 266.986244401803, 
    265.212200603685, 266.493623591346, 272.288149829089, 273.386152478814, 
    268.924946560023, 266.18827640176, 263.691989549393, 266.285618930293, 
    272.147235596241, 273.128562047982, 273.28560958424, 268.877592318825, 
    264.122921704056, 265.451751740062, 270.262857290283, 270.394338439117, 
    268.445325138126, 270.343877817861, 263.923905131508, 259.724714569852, 
    263.410302497811, 265.145636140635, 267.903671741883, 271.444698693992, 
    268.796101741652, 267.272988715779, 266.671097328722, 265.857691771694, 
    264.696211018142, 262.441452462356, 265.995678086382, 270.697580559426, 
    273.548544348543, 272.335679816075, 268.082412864782, 264.833791787064, 
    263.931991736281, 263.493322186025, 265.619303139004, 269.153551721494, 
    270.255766279264, 270.635853683275, 268.546794508335, 264.468344533033, 
    262.094398287137, 263.188995274788, 262.678016991877, 261.590956645405, 
    262.601978156707, 262.831407650722, 264.127196888447, 266.687009171795, 
    266.203775066216, 265.810355496317, 265.235557340887, 265.616658478407,
  256.476329399155, 263.189577026059, 267.286601984013, 268.148857942004, 
    267.819463510873, 268.2964470421, 268.891061935158, 267.270860822703, 
    263.880282948851, 262.357727244434, 263.895338186966, 267.720010477863, 
    269.176185329385, 270.182413483618, 267.692981560128, 263.972755111048, 
    261.265059164556, 261.326433981209, 263.213133216403, 262.992297948421, 
    265.209087437873, 265.042465570897, 260.980010052506, 260.996270496626, 
    262.846168210395, 264.720072782916, 268.2186758597, 266.510298656241, 
    264.986835190787, 264.505334206333, 262.520721327345, 262.088153095239, 
    264.088389016534, 265.44880297916, 266.834086170022, 268.001125821257, 
    268.248644571196, 264.274737881605, 259.859581372858, 258.947436860164, 
    261.437812035252, 264.118736957055, 266.350333530163, 268.452789996646, 
    268.047883068697, 265.654800170958, 262.685195508205, 260.476694828711, 
    260.770408473498, 260.95795550415, 259.055488258207, 258.883048382092, 
    259.442145652713, 261.041772920786, 262.569936007053, 264.118868614028, 
    265.21496703119, 264.60288828208, 261.940583284178, 258.600625378939,
  262.459304103509, 263.641709172015, 264.981954273331, 264.705423714311, 
    263.812371032295, 263.57534769206, 262.357752737938, 260.148951731588, 
    260.711967688372, 262.344123198653, 263.133182032455, 263.85789596085, 
    263.405724854136, 262.72330566662, 260.020591441197, 258.650555374814, 
    257.637752648132, 257.241765658466, 257.76330400005, 260.00914142633, 
    258.460561053046, 256.865072147695, 261.577524848764, 264.012413037364, 
    264.419737837483, 264.871199612601, 263.872378074493, 261.701176096106, 
    261.819563754279, 259.811408945657, 259.687231925287, 260.021452135096, 
    259.740028112614, 260.374336702377, 260.469535381265, 259.107602756199, 
    257.149745119566, 254.812167894857, 255.376365003159, 259.320083808014, 
    262.461337583191, 264.498309240072, 265.277349656251, 266.083346425238, 
    264.313022735939, 261.151727556101, 258.535421011435, 259.491117642337, 
    265.721448196726, 267.030928180724, 262.803914643381, 263.73265805612, 
    263.164385746492, 262.935211696302, 262.974553131615, 262.395900669062, 
    262.288264400873, 261.315773281852, 260.409792978253, 260.913455394112,
  259.577984950304, 260.7278246248, 262.134847104423, 261.064398415997, 
    259.693379621545, 259.02560487763, 258.29292838359, 259.056655424913, 
    260.679460786829, 261.44059636255, 261.574107459471, 261.163089737056, 
    260.424400737215, 259.304937325989, 257.318268336393, 255.447576811254, 
    253.805248981622, 253.330192731882, 255.27066780075, 258.935278747472, 
    261.049683545994, 261.250509469791, 261.84005936589, 261.770395161248, 
    261.360954107844, 260.437717144241, 259.319853228964, 258.320725771499, 
    258.170597984571, 258.111275264748, 258.491288390506, 258.448510532413, 
    259.254327832421, 259.913589211694, 257.804264000891, 256.248817814755, 
    254.043262173108, 252.280318013137, 253.917667128914, 257.319981305811, 
    260.836673545457, 262.727187596796, 262.528268509599, 261.529818949403, 
    259.458402434794, 258.161870778386, 259.616727935719, 262.864345251921, 
    262.685110104377, 264.678991489571, 261.587871835912, 259.773676788833, 
    260.766099438121, 260.942179044089, 259.837978011666, 258.609175817479, 
    259.179541014736, 259.568749365777, 258.683844572258, 257.644924314444,
  258.064427100439, 258.925439949305, 260.123371740646, 258.749991249001, 
    257.123993679831, 255.797704919887, 253.697499928584, 253.594832296819, 
    255.969709008359, 258.345576575168, 259.715238256689, 259.54889698447, 
    258.66512437667, 257.500036526207, 255.906551013681, 254.753608560064, 
    254.877309856316, 255.282151671368, 256.485774539163, 257.858984266652, 
    259.171272111867, 259.261949127642, 258.768366983477, 258.577919692285, 
    257.574823202309, 256.999750216431, 256.439030534162, 255.580433291305, 
    254.913671419411, 254.574396732796, 254.867302348775, 255.502984831696, 
    255.258217767699, 255.063684734503, 255.787847943009, 255.861369585844, 
    253.151678124325, 254.793103843154, 258.213765313787, 260.129503423322, 
    262.814060267515, 261.87663069152, 262.41574994121, 263.254376413115, 
    262.104055334926, 259.745359300549, 257.779461235934, 257.653846950031, 
    259.26060983541, 260.409029215129, 258.9594488671, 256.534434000958, 
    254.866675696098, 255.189389648836, 255.546993782339, 255.693384923203, 
    254.780976203783, 253.999495305391, 254.351191991627, 255.363400081092,
  252.342273816056, 253.629429407269, 255.215355340308, 256.149376061891, 
    255.855482989067, 253.717695330484, 250.277986256936, 248.502430543001, 
    248.609569959765, 250.385300082035, 252.767090845517, 254.664462332567, 
    256.042869268451, 256.713154602749, 256.580238175941, 255.469183334059, 
    254.962617352347, 256.323439358937, 257.845299796446, 258.562664861725, 
    259.240365951142, 258.72414520324, 257.790015503492, 258.156370717706, 
    258.803404343178, 258.95553808949, 258.360186911814, 257.21342136238, 
    255.730826020227, 254.322250570323, 253.360715234451, 251.850028668112, 
    250.028441999848, 250.730394623364, 253.392045224801, 254.417320494165, 
    252.007806995298, 249.438691217469, 250.109681789122, 255.619085676633, 
    259.440640009618, 260.464430366332, 261.711557391732, 262.471163769669, 
    261.495020480976, 261.235926508626, 259.946753741146, 257.846788083662, 
    255.997653042129, 256.023319650562, 254.934721441523, 253.101810707019, 
    251.418161104608, 251.097469734341, 251.016007938658, 250.058857437973, 
    248.857744276231, 248.054796031198, 248.560375718746, 249.891595417045,
  248.729010292848, 249.00229060877, 249.688401308299, 250.462800214652, 
    250.545027035681, 249.938828370831, 249.446525284193, 248.594661210062, 
    247.074944961913, 246.496463235658, 247.356944562831, 248.632223697731, 
    249.725465970968, 250.3239432273, 250.020884908765, 249.125859239913, 
    249.310762131669, 250.243700462585, 252.423988921495, 253.975950982616, 
    255.259222150423, 256.259499927434, 256.643262029456, 256.788826837781, 
    257.046242335316, 257.084371447719, 256.668006907982, 255.993719772485, 
    255.627301064576, 254.534839950128, 252.892377872552, 251.364768639366, 
    250.196408375235, 249.839306017373, 250.380833985085, 251.135462130128, 
    251.003264720371, 251.161618758164, 250.650889811433, 249.437722307561, 
    250.144785391273, 251.739337869848, 252.696554126473, 253.083090956952, 
    252.888630055344, 252.415539112652, 251.630686028373, 251.640230362371, 
    251.998378264956, 252.364844260499, 252.314302376377, 252.830895892491, 
    253.349171992794, 253.256328517409, 252.680821544148, 251.696783696199, 
    251.716080090265, 252.037659250574, 250.277410970508, 248.578026632474,
  248.060913425689, 247.205823554775, 246.925430023324, 246.855186690582, 
    246.906628258783, 247.119728927982, 247.521560689479, 247.943244836837, 
    248.41072010727, 248.671774967141, 248.621110147825, 248.680055137634, 
    249.052212825149, 249.531294519588, 249.948619425968, 250.300511404811, 
    250.573455756581, 250.448254602621, 250.562173695695, 251.072371059435, 
    251.754008281051, 252.521162992005, 253.092794605794, 253.49704162634, 
    253.580585286827, 253.51825998504, 253.378768952599, 252.595846363368, 
    250.736279883955, 248.866608888955, 247.794709443619, 247.172428984507, 
    246.604329423242, 246.235499508915, 246.168888743745, 246.342045799954, 
    246.7813764648, 247.691682348288, 248.620079318172, 249.115694874972, 
    249.075755768763, 248.804852423344, 248.857589245107, 249.251081164037, 
    249.646479135133, 249.956603690843, 250.074078268057, 250.088368656717, 
    249.935008035755, 250.04478851018, 250.571763211736, 250.991117817773, 
    251.143954031713, 251.224230649496, 251.031393799222, 250.647806154737, 
    251.342200483882, 252.8825666317, 252.438370392729, 249.963057567157,
  247.963796648906, 248.596038865446, 248.750001169468, 248.492097204227, 
    248.303646072946, 248.147733339006, 247.90722353499, 247.729796184756, 
    247.731094263983, 247.77310518122, 247.707258758209, 247.508382074215, 
    247.354119112971, 247.284994415045, 247.240760970344, 247.18649599188, 
    247.151004618765, 247.062688695634, 247.053188908177, 247.22091541464, 
    247.450229257327, 247.661044761903, 247.833932568375, 247.884154752323, 
    247.874827656156, 247.707312520157, 247.324885674037, 246.730502986875, 
    246.324280932454, 246.316255943322, 246.806820493277, 247.409612414815, 
    247.722156352814, 247.663286680425, 247.484906960977, 247.401463855404, 
    247.482355505624, 247.645021782041, 247.787470104492, 247.784938548059, 
    247.651692447999, 247.508737033241, 247.489772830068, 247.455501521042, 
    247.436620417439, 247.477650480924, 247.505128421651, 247.508325848573, 
    247.451568196191, 247.480426131897, 247.520336724811, 247.588910730406, 
    247.840031643419, 248.077666696089, 248.276980306636, 248.473979333648, 
    248.690377684765, 248.496174920054, 247.877844737354, 247.562253644704,
  259.652698229391, 259.686423991075, 259.749603034073, 259.768963031064, 
    259.736418532164, 259.620753596576, 259.501736493651, 259.229485323511, 
    258.922992359888, 258.652642221336, 258.448444235645, 258.191451502576, 
    257.968267899341, 257.748822330411, 257.580066815981, 257.709231414371, 
    257.679883806486, 257.775162577388, 258.421296179659, 258.864474209832, 
    258.426337482306, 257.939188764022, 257.706461131264, 257.843076044175, 
    258.208907237615, 258.623200573519, 258.926165272898, 259.094551735915, 
    259.120654577766, 258.765207766704, 258.178908974232, 257.617496110077, 
    257.148015206318, 257.138846529594, 257.578441941942, 257.81955048862, 
    257.879272852889, 257.823613726265, 257.797389891807, 257.70915755931, 
    257.607894361407, 257.465557268162, 257.389109220489, 257.359135401235, 
    257.405799895267, 257.376162352535, 257.289848808647, 257.249547155327, 
    257.357413576945, 257.554177115258, 257.756938652061, 258.015639904705, 
    258.278050759179, 258.523331876126, 258.783621134737, 258.996598794731, 
    259.185049344684, 259.388082848557, 259.534564599326, 259.621092875782,
  262.804884193871, 262.365493541927, 261.654113932089, 261.213746265513, 
    261.142958502872, 261.421021665638, 261.477016164053, 261.239749542805, 
    260.51798714719, 259.539460215319, 258.898605149899, 258.622629712321, 
    258.558449119521, 258.75514226013, 259.103529130753, 259.802112061606, 
    259.874053867642, 259.344117618246, 258.38137047264, 258.285446737498, 
    258.592608225664, 257.326674517145, 256.319642629491, 256.561488735162, 
    257.278848214193, 257.720481851729, 257.62898034324, 257.309407425171, 
    257.253538817783, 257.379142517373, 257.570943710091, 257.946412646657, 
    258.090117620254, 258.310997756774, 258.951304738272, 259.525531238296, 
    259.840744446095, 260.134672308369, 260.721729973691, 261.134809168288, 
    261.423267624934, 261.54358767906, 261.598668997779, 261.762202283977, 
    262.265853897327, 262.826599518545, 262.992407673186, 262.897289680089, 
    262.816378275645, 262.756311348635, 262.680742015355, 262.599276582176, 
    262.637562240319, 262.779355436532, 262.841961137808, 262.941653793907, 
    263.018813491984, 263.024880025055, 262.939894975731, 262.889110410311,
  265.346641410352, 266.98331766661, 266.616146355981, 264.958067941705, 
    263.729777170238, 263.808298016044, 263.731410954181, 263.102626975933, 
    261.100554277546, 259.006296386024, 260.601090345654, 262.507746711193, 
    263.250459871422, 263.140022280079, 263.419707277603, 263.372963209835, 
    262.663227300322, 259.760501914299, 252.163416967601, 255.172765460205, 
    262.361609035064, 261.170558020819, 260.917205319054, 261.674619465723, 
    261.781725878668, 260.999939446314, 259.665419732649, 258.346622146717, 
    257.587898718319, 257.542083910435, 258.378331007823, 259.175552766469, 
    259.824431614896, 260.100386154124, 260.24717314722, 260.556538947079, 
    261.074029797192, 260.605918754215, 261.385962893625, 262.918194248748, 
    264.075318958481, 264.362813575888, 264.075078671532, 262.974136916087, 
    262.489226837092, 262.709264923131, 261.734561715911, 260.998490083758, 
    261.328476047796, 261.198093444113, 260.792936488475, 260.377179908775, 
    260.073472993599, 261.612038410479, 263.095777562588, 263.350995354205, 
    264.930482401901, 265.68611142123, 264.507231053127, 263.877622725058,
  265.306747718412, 264.696930862651, 265.211844580424, 265.893939647171, 
    265.106099905033, 264.750431634797, 262.134670294383, 259.952030256444, 
    262.305422268417, 269.012416233867, 270.85178672414, 268.128483928344, 
    267.605012173643, 265.124432491104, 265.126349735778, 261.964308132941, 
    258.042309430409, 262.120089506995, 265.346695111987, 269.032432334489, 
    272.866393530019, 271.218645589967, 270.440564368522, 268.448590799549, 
    267.609373598005, 266.242716327301, 263.994232220326, 263.385532611277, 
    261.203045730303, 257.709305839886, 258.226208418137, 259.490401097355, 
    260.137247759042, 259.91320014223, 258.853678084371, 258.342020081322, 
    259.68207106502, 259.621680188893, 262.583413607305, 266.695801215618, 
    267.838438342766, 267.584759795841, 267.475564717332, 266.0832822405, 
    263.434853810177, 262.702241065079, 264.514276911803, 266.020193705241, 
    264.401808999733, 261.236462838027, 262.610719982996, 266.392351202465, 
    267.519219578794, 268.772221926496, 269.083837005907, 267.66860859753, 
    267.564598297408, 264.584077577813, 264.06031474945, 265.525657720017,
  268.817382960363, 267.969660300008, 268.181629172648, 267.594207266302, 
    265.058399357766, 262.00217512344, 260.280496462267, 262.107281372674, 
    268.113027190393, 272.847867663063, 272.138394630096, 272.476783770124, 
    269.212279165256, 264.604258350839, 264.980595088977, 263.609447052339, 
    263.431681165748, 268.941541639647, 270.521527841469, 272.627179750263, 
    274.947596032549, 274.780463010417, 274.395335524046, 274.346247662081, 
    271.842638886238, 269.346798317772, 270.234498456755, 268.98635895911, 
    263.640156060843, 256.715162649777, 256.238087206505, 260.1013061214, 
    261.158170548514, 261.355333586198, 261.338599270632, 260.995054878012, 
    261.936426765434, 264.972351884475, 267.81839587252, 269.409530734619, 
    268.476893301459, 266.996436548416, 266.698768759536, 266.013006834871, 
    264.795770198046, 264.742581439496, 265.178682603665, 265.070449081445, 
    265.750338580617, 267.995649485192, 271.271472516825, 272.127684473452, 
    271.118280106129, 271.829163973855, 272.565717947145, 267.272486635743, 
    265.67051278109, 269.195507358241, 270.463210334274, 269.748593010421,
  268.632667111825, 266.86396032502, 264.460797686824, 262.744416863158, 
    262.372256967353, 261.850578927627, 262.216693993989, 263.812862090047, 
    271.797468167939, 277.428251182839, 277.619195384865, 277.515807972056, 
    273.610804205372, 268.040543269307, 265.640573392647, 267.381793491711, 
    267.658076481985, 271.364108792855, 272.221810740941, 273.747845776335, 
    274.872842489737, 273.111966628293, 270.556577188632, 270.11775285153, 
    270.757170685111, 271.839941153082, 274.225030852854, 266.310766312396, 
    259.919610906891, 262.471618096464, 265.677560395468, 267.639894816477, 
    268.10381033241, 267.621557588165, 266.611457406597, 266.818660067887, 
    266.768632304769, 267.999293428557, 269.337746023919, 269.460124796381, 
    268.294697113616, 266.740431595778, 265.459317918515, 264.821377588259, 
    264.627435404849, 265.297672822921, 266.124983972916, 266.787149511768, 
    267.425178140729, 269.171389049837, 272.351586381717, 272.116359017423, 
    270.726713395509, 268.837219473499, 268.307576118762, 268.576798222416, 
    270.385384546411, 271.436526858654, 271.276153864959, 268.826814952394,
  270.417016119965, 269.571760154537, 266.823345525021, 267.429094950204, 
    266.578917276757, 267.406172198589, 266.789120432033, 264.916276243501, 
    268.905352502367, 275.94349907601, 279.047740813467, 279.74597788761, 
    279.044305448572, 271.997992064778, 266.371871589955, 267.462959399603, 
    268.612761958002, 273.383529769305, 273.654890202308, 277.049750760475, 
    275.998738542689, 274.321814169672, 270.499670971558, 269.536384716154, 
    270.51305482187, 268.255885289963, 265.60460675834, 261.585921181245, 
    262.186090063168, 266.829938478814, 270.974534084908, 270.986952335243, 
    270.136942496485, 269.045267566917, 267.328464236061, 267.583129123503, 
    267.938193359658, 269.758008858711, 271.165669079076, 271.085642605941, 
    270.68811563868, 269.081360926102, 267.00262616609, 266.486449670059, 
    267.240650594629, 269.43124714966, 271.23147383283, 272.221309133956, 
    272.186333369896, 271.179004149532, 272.980784436945, 273.405496507433, 
    272.043216985559, 269.97272040623, 266.409355922306, 268.987105008573, 
    269.821234182646, 271.792343162243, 271.943626046032, 269.780056590371,
  280.006001343351, 279.397263136418, 273.4672409874, 270.823214198145, 
    269.802296773484, 272.866723455767, 273.611556970151, 272.849363489424, 
    271.63748486117, 272.056910487831, 276.221664730406, 278.966906971021, 
    275.495744039294, 280.215865556628, 276.30488211079, 268.839063910806, 
    268.325414364849, 270.431332048533, 274.123573992315, 280.594606403997, 
    279.265134661551, 278.394061095522, 275.979832451571, 270.669461367684, 
    267.031597313925, 264.295651428531, 263.823217767752, 263.336798093962, 
    265.353351807346, 270.478257056065, 275.204657648402, 275.032084658683, 
    273.087380764749, 272.833958257287, 271.781913521658, 271.689876575121, 
    271.837272724874, 271.939822742534, 272.861594429022, 275.789349197436, 
    278.404642345512, 277.054188981033, 274.14227644506, 273.601571344397, 
    274.962232454542, 277.233180322967, 279.285576135351, 279.979544154802, 
    279.602984939643, 275.790684089798, 275.323077824468, 273.278160486913, 
    278.578540964102, 277.320222737842, 273.696550580148, 270.718731940866, 
    268.632731170482, 268.359174158345, 267.208739113815, 270.88476131248,
  280.006116812236, 281.822748003017, 278.580581224384, 277.693022452066, 
    278.906304682158, 279.885643751047, 280.035093818202, 281.570791558376, 
    278.158573566384, 274.555084407326, 275.781277072891, 280.893808049529, 
    280.2075009779, 277.412364734971, 281.580380041718, 280.540448983047, 
    274.708796019788, 274.357893093645, 270.097673925208, 270.445784790379, 
    270.58442953352, 273.621069595859, 283.079433033547, 280.546413340593, 
    272.445252310679, 269.770640492707, 272.039614686014, 272.95337995766, 
    276.442475969428, 278.666617060412, 275.875073138039, 278.49535756583, 
    283.557558796989, 283.699862749083, 281.37382794477, 280.642682083671, 
    281.136990106979, 279.367733859381, 276.213341137201, 275.000202181744, 
    277.098068024394, 280.582613866415, 281.893080010947, 280.48643751426, 
    280.400768250201, 280.168192494159, 280.522590864364, 281.983761571217, 
    286.698768830106, 284.995443013879, 279.56382645303, 273.554929748303, 
    276.609605194066, 286.109162808372, 290.127508743395, 281.955367693257, 
    277.985356790229, 272.020388404432, 268.213207107958, 271.080016775142,
  288.698573820288, 290.17547871823, 284.591253388761, 282.445356877165, 
    282.932453507582, 282.47855901466, 284.607563127178, 286.895670834222, 
    286.32180466823, 286.155599470804, 285.697588619111, 282.116860304239, 
    278.556002271479, 277.128042138512, 285.638481733707, 290.192587073433, 
    284.226209918631, 275.414497237197, 272.095744706789, 275.708905025306, 
    271.553958625837, 271.426196640184, 279.646076061455, 284.555239820046, 
    283.017285553636, 277.377741213537, 279.246748516478, 284.240730571531, 
    291.160127857579, 293.785820796848, 284.247138889185, 275.600950567513, 
    279.401323699188, 282.528908088769, 277.823591929023, 279.740743741994, 
    288.989599786444, 289.02174827416, 284.064017285557, 281.431808190949, 
    283.688053294607, 288.788738863842, 289.714645297116, 285.373293694126, 
    279.701233329003, 278.489103291319, 283.753779892985, 281.950453965805, 
    279.117515686457, 285.835837942949, 286.075750227435, 281.566480894604, 
    281.371811325028, 289.570110819461, 292.760474382914, 293.250063073564, 
    286.430815615811, 277.77245858377, 274.208087316662, 279.212736049695,
  293.933658259651, 293.672893082636, 287.519268204053, 285.970700798461, 
    289.198512683594, 290.789531039818, 290.823688448131, 290.419134582231, 
    292.505688663699, 292.831610288311, 285.821011174558, 284.458656958837, 
    286.014055023219, 286.224007716923, 291.415868336935, 292.193919291432, 
    289.306250322175, 282.033296158576, 273.937733670164, 271.331770346385, 
    283.945870564824, 292.445364205907, 291.258424761784, 288.327020619715, 
    286.976071395065, 284.760526306352, 280.209239937356, 283.51060878638, 
    289.35291510295, 294.398290146938, 293.478779852946, 286.11040280555, 
    285.899373393355, 283.799738409756, 286.187267692081, 290.595636531669, 
    292.963010417126, 291.011685350898, 287.001736178611, 284.972764246443, 
    287.110248533294, 291.490810138468, 293.641936068103, 290.658134475034, 
    286.59923069714, 285.086313522099, 284.2846314565, 286.014876127163, 
    288.001995132156, 290.987114077999, 290.008904820435, 285.653030379881, 
    283.574468952549, 289.368758730261, 294.505442558516, 292.72471647515, 
    289.873069411844, 283.969839822372, 281.097302481738, 285.401387141191,
  295.226249374011, 296.032094878916, 294.599832741624, 292.378995106991, 
    293.602634504489, 294.629651454567, 294.187191955438, 293.692020652679, 
    293.483101152949, 290.795489453025, 287.735465912344, 293.100616994658, 
    294.54748778418, 294.605851986711, 295.317913628682, 293.464020080107, 
    290.129667107867, 285.086483361337, 280.271251861898, 287.264155071818, 
    295.194808544435, 291.177348510701, 291.216466852779, 291.083590034377, 
    287.866091432673, 281.091620490657, 282.613106656032, 294.796566967335, 
    297.758783628323, 294.26469809539, 295.136409535843, 293.095891737464, 
    289.945407402595, 289.200157197819, 294.830301823264, 296.874483964825, 
    295.198263524997, 295.14536462865, 293.183199230001, 292.388932198323, 
    292.338340263186, 293.384318652065, 294.403644128336, 294.277776579418, 
    292.073600855593, 289.720303113853, 291.132685770923, 294.074450062181, 
    293.446795387289, 293.536698347528, 294.491552614406, 290.140965038041, 
    288.741762462986, 295.086400761671, 297.445736099515, 297.365993668628, 
    295.071035821556, 290.193118457963, 289.58857319414, 292.008739526228,
  300.378562114835, 298.628901774598, 298.274301595821, 297.12445438714, 
    296.637140296089, 296.549929531784, 294.454056405968, 292.214680021402, 
    292.411415697051, 288.458906797274, 291.489151355905, 299.685799917374, 
    298.946922708895, 297.35479621966, 296.655249245296, 296.056811190784, 
    292.399195445851, 287.80530244723, 288.961947582226, 299.421924886053, 
    297.99865239338, 291.395759957297, 291.410553936795, 292.348669332452, 
    286.799630374231, 283.783430084043, 293.767236581966, 299.98156008976, 
    300.792457385189, 296.955699379386, 294.845197343338, 293.498402962016, 
    292.859064383138, 297.346266774055, 301.775150076595, 301.134807965063, 
    299.487819310837, 298.457234121202, 297.453354227585, 296.48430697036, 
    297.838755113959, 298.602992743257, 297.447812377709, 295.440665770367, 
    294.022242743605, 294.901845753064, 298.515928915959, 299.984462934551, 
    297.628982064338, 296.285417716879, 295.631573552532, 292.923771557041, 
    295.86944632705, 300.799445771948, 301.079087599678, 299.597850020762, 
    298.090412004476, 295.400493408451, 296.138569097958, 296.234253752241,
  304.533475117741, 302.15133996765, 300.427900766823, 298.893111175541, 
    296.698214490675, 294.564171428032, 295.227257207017, 294.956627119894, 
    293.488435206752, 295.566600689206, 301.394316839548, 301.140142826778, 
    298.80608276937, 297.524705578044, 296.174191168213, 295.366920931531, 
    295.091711513046, 295.515389745006, 299.82680398518, 302.086350687554, 
    301.899333423735, 299.346208509808, 292.871157175425, 295.144387937969, 
    293.113835792816, 298.01162652582, 303.213445237065, 301.645064103065, 
    301.260106656916, 298.390076569884, 298.05979261671, 299.21185146887, 
    300.917595902536, 302.192307851227, 301.287328719171, 300.678334810365, 
    300.669297146292, 301.058456248634, 300.827208936125, 299.749546796703, 
    302.04261396018, 301.616395902016, 300.938737029755, 300.297990434174, 
    299.69369238642, 300.990825678062, 301.416203022972, 300.187663435738, 
    298.773713647136, 299.127423610331, 299.153996909499, 297.737288417111, 
    301.556802731031, 303.818712227912, 301.922469874234, 300.718497377957, 
    300.26466559701, 299.540641596708, 300.346686033526, 300.346734194289,
  304.000122460167, 302.832245895577, 301.490970250057, 299.996748729579, 
    296.974901303133, 299.183457441297, 301.486243870238, 299.251876033658, 
    300.055149566375, 300.504151294353, 303.582404793059, 302.758907736999, 
    301.522053222464, 300.658551516823, 299.741812196675, 300.200717110373, 
    300.164583826671, 301.103522258481, 304.538807852741, 304.773227743231, 
    302.858134398201, 301.023353205772, 300.09422004086, 301.73886252402, 
    301.431019322744, 304.014692512592, 304.267379896907, 303.842320834391, 
    303.142127314918, 301.921333939023, 302.093870553862, 302.857812697288, 
    304.641815494924, 305.179996895878, 304.1965496882, 303.367147037545, 
    303.377404401283, 303.819614537244, 303.267886671206, 302.742978437826, 
    303.016943294174, 303.24977993837, 304.417873443292, 304.123187103624, 
    303.709207405139, 304.898409204226, 304.239244265843, 303.262793490016, 
    302.890701647178, 303.297209447782, 302.92381423827, 302.035255482978, 
    303.660466476532, 305.664656099911, 304.443935242904, 303.74054992196, 
    304.020751819188, 303.996832497205, 303.473541745381, 303.578003739516,
  303.005590048383, 303.932360520834, 303.315660968529, 302.082048776738, 
    301.832415090835, 303.260485354026, 302.549105378987, 301.204946840385, 
    300.071747928248, 300.135831899164, 304.047382109009, 304.636960789334, 
    303.957513746329, 303.600641879097, 303.469728601454, 303.240278685217, 
    303.593412300415, 303.529048083934, 304.40453014428, 303.867298347714, 
    304.53775862636, 303.282202103877, 302.929322269922, 304.82962726739, 
    304.52589865887, 303.97873118273, 302.63904288696, 302.438303518401, 
    301.910142356216, 300.862922211985, 300.531770956833, 301.144096280433, 
    302.882147214886, 303.9803877411, 303.7882124389, 303.660478864527, 
    304.185393298779, 304.210924796954, 305.496073017343, 304.463722139271, 
    303.418637393892, 303.484666025835, 304.828382083749, 304.410380628051, 
    302.802077143627, 303.274403240799, 304.17357567133, 304.125024536135, 
    304.060786873019, 304.099880871655, 304.33771001193, 303.973891628247, 
    304.429325359796, 305.111233221674, 304.495574570154, 304.391250701577, 
    304.462085005271, 304.264184865012, 303.429872173247, 302.820017569888,
  300.630267118268, 296.530815263696, 302.421111039314, 302.034325489507, 
    301.929992498916, 301.986241169021, 301.07464869478, 301.855029042397, 
    300.556019634788, 301.424884782174, 302.59897156449, 302.651175476358, 
    301.678908408495, 301.060904677731, 302.013154444408, 303.048057199135, 
    303.002082839862, 302.275032392774, 302.498481082659, 301.620614546937, 
    302.277602479178, 300.592643539355, 300.625629427117, 301.956091729326, 
    302.252117031072, 302.226134587006, 299.033484302033, 297.88258828675, 
    297.659958107026, 296.433806450229, 294.823669370521, 294.290033259598, 
    300.483159188289, 302.347585782199, 301.668717013895, 301.388968198182, 
    301.762731798883, 301.175102125952, 302.166640493609, 301.796217104552, 
    300.947335458338, 300.474529248065, 301.943427486891, 302.071116722553, 
    299.988578000387, 299.600721102289, 299.847949720793, 300.686139246326, 
    301.546790907126, 301.71603525185, 302.762449143469, 303.028287955578, 
    301.645153735198, 301.189556258527, 301.761753728422, 301.783313157281, 
    302.117018034919, 302.77657146901, 302.846624767307, 301.33420919893,
  296.474261618152, 288.807071576618, 294.757199386662, 298.024123899055, 
    299.355393391733, 298.602270031105, 296.701749716705, 295.381788258869, 
    293.048261416428, 293.215652076, 297.661371762091, 299.090528471803, 
    298.377054120538, 296.445544488254, 297.586691769479, 299.85843013531, 
    300.288518060003, 299.765695860969, 299.373235854293, 297.82346741776, 
    297.497978397216, 296.794902393392, 296.64582025307, 297.757826421303, 
    299.503222794413, 299.404353429061, 295.881960055771, 293.862623843874, 
    292.303030565755, 290.369812467162, 288.69275808675, 286.748029690007, 
    291.466454206, 300.027067471447, 301.106732406375, 299.41560230197, 
    298.851119968504, 297.503056358463, 296.525617119111, 296.340996819052, 
    297.234644500508, 296.82315778787, 297.785162633995, 297.576777748732, 
    296.042833079314, 296.014090992179, 295.518115038767, 295.764160754625, 
    297.22165264933, 298.808068975035, 299.726406912336, 299.367226347577, 
    297.070944322677, 296.557026270671, 296.35664702987, 295.634384082233, 
    296.49599924064, 298.418820340937, 298.206385984131, 297.112902636801,
  290.057827883747, 289.218290959649, 286.807164889107, 288.008063570125, 
    293.671614256244, 294.503927928323, 291.21176563549, 288.427885108786, 
    284.875513786345, 281.69518448895, 286.102628295131, 295.278029735836, 
    297.532078400881, 294.849515188796, 293.105275248942, 293.151250873541, 
    293.346730029769, 295.664490048899, 296.481553976194, 294.535443981384, 
    292.932132318515, 292.04714793346, 291.588456498433, 292.582106332476, 
    294.508268793452, 294.848638872323, 294.236217306917, 294.221892508247, 
    291.269117126872, 288.420587520874, 286.017099605289, 283.745831782976, 
    282.254537380486, 290.471229633952, 296.97637913093, 299.120285503912, 
    299.542721850048, 297.744549263445, 293.811798043652, 290.269477059666, 
    290.448406670928, 292.358735570612, 294.348801798082, 294.789914424452, 
    293.746124688521, 292.524029024049, 291.721970521648, 290.386678748769, 
    290.811962800316, 292.152841550995, 291.334743097911, 292.147317762903, 
    293.65561389907, 292.94601113018, 292.574635811808, 292.379754362886, 
    291.866651490783, 290.549448037314, 291.724901061077, 291.678817482587,
  294.151843894314, 284.538948166965, 279.248852183482, 278.423333356182, 
    288.425322488314, 291.664434977229, 287.587950391837, 286.302235132601, 
    284.61681297687, 279.183529181634, 276.466271286113, 286.893094541808, 
    292.619788682365, 292.230290550611, 288.385283011625, 286.231771312061, 
    284.708906070485, 287.785155567552, 292.974918240042, 289.502744269138, 
    286.029122414765, 283.301524146869, 280.78609609719, 282.731446217734, 
    287.986569586195, 289.047197523121, 288.253187944906, 291.439177202533, 
    292.573855592884, 289.75845166343, 285.215906118637, 282.908575944042, 
    279.281628386521, 280.462078477014, 288.052015208894, 295.188158548048, 
    297.981207325464, 296.137253270621, 291.874160610095, 286.627017301745, 
    282.616854158787, 284.239789953386, 288.737151174122, 292.985891743519, 
    293.740606970691, 291.206676106466, 289.796790712288, 286.145384488586, 
    283.00405638528, 281.705718405608, 280.779144764431, 278.618619562509, 
    288.552730885287, 293.315636379319, 292.082383152576, 290.658504678513, 
    291.951233514516, 290.22107459677, 281.286509862024, 288.92964215283,
  281.103090422496, 272.176049218727, 277.693934997084, 276.121419441018, 
    274.134695847777, 282.081211226202, 284.906131115347, 285.888758448112, 
    283.019850010895, 279.054878686578, 275.643992826325, 281.208316927457, 
    290.329850015604, 286.845410802421, 281.140146689295, 280.528062188574, 
    279.848841825509, 275.623507353461, 281.8072153939, 286.431969773206, 
    281.253711161875, 275.672804890889, 271.867775170165, 269.215051651129, 
    277.256072895995, 281.964197235466, 282.551907111959, 287.170957583914, 
    291.817169683166, 287.66302078205, 283.680589059478, 281.743932011296, 
    279.015473550084, 276.570468419745, 280.525827714384, 290.292197576631, 
    290.905317837906, 286.607656522541, 282.638998027849, 283.044069707496, 
    281.587213462674, 276.894898825205, 280.517115423544, 288.802956208227, 
    287.691276142715, 286.510768496536, 288.943646621373, 287.973320221018, 
    280.435875440815, 276.366182955841, 273.473280156091, 266.141072729037, 
    274.166520744228, 284.261350782433, 284.810197821948, 286.520963891097, 
    284.445547364948, 284.412737782882, 284.579115724753, 286.338674342218,
  271.565234762739, 272.332890068602, 275.60412701381, 275.146663911133, 
    269.078852379109, 275.624176686704, 285.127092032282, 281.980660210745, 
    276.320102533934, 275.20752924475, 278.904465942612, 280.760831915058, 
    287.484670814855, 287.795643853211, 284.002941709951, 277.333180377561, 
    275.091946538885, 278.264779442277, 284.45875912297, 287.322079567602, 
    278.889454189652, 273.059558803857, 269.562196632915, 266.181588416897, 
    268.491683548257, 276.951629304431, 280.242971577324, 282.964166111212, 
    281.809607904099, 277.483352515044, 278.515881853163, 276.697174890997, 
    275.279279949516, 277.475611003929, 284.213673595049, 288.212607370318, 
    286.202703014318, 282.227345357384, 276.043782507941, 274.693287415442, 
    275.53126556803, 271.629811174734, 278.333787961057, 281.872820709192, 
    286.739086779711, 283.893573224656, 276.448043290263, 274.95380329328, 
    272.748713491889, 270.415448208984, 269.637041922257, 271.076140868905, 
    272.461953525318, 269.157689511333, 274.224911541735, 279.149804624438, 
    273.825390221774, 273.917406046507, 273.046670647437, 276.262723839094,
  267.825686085268, 275.989279342754, 280.824385103457, 279.291215250768, 
    278.373195161016, 278.447399027565, 276.709094691406, 273.293807134234, 
    271.896996252893, 273.056598583974, 279.63006840689, 283.751047314292, 
    283.382631625205, 279.63353796934, 275.994752291691, 268.730049115037, 
    265.533835245261, 270.186093281154, 275.326984658625, 277.524732196334, 
    277.673883512546, 274.584884630725, 270.763884271627, 275.69489755256, 
    276.862386741293, 276.580308510986, 278.803587665789, 278.923623017741, 
    273.756545671812, 274.583255251978, 274.542812111094, 274.576311538128, 
    278.215427446816, 277.927853520426, 278.309818340325, 277.227144536833, 
    274.240993308284, 270.496699985122, 267.84150558872, 267.33614520097, 
    271.585943200867, 272.313554106014, 279.161735283571, 285.851436940304, 
    283.188766716254, 272.298134874434, 270.203850718307, 267.070200706542, 
    269.801280577925, 269.858826519894, 270.730871774505, 272.500067459896, 
    271.112670367704, 269.506115435182, 275.052156971377, 274.164360893186, 
    271.912879504993, 273.098008780213, 268.57159111665, 267.824712758921,
  268.364303705136, 271.563020097995, 272.65346950918, 271.950467165418, 
    272.154984610938, 270.377425145637, 270.208931577868, 270.548932093834, 
    273.441870159344, 272.728349702, 271.571044994246, 273.282461255919, 
    272.600958760403, 270.263036706784, 269.621896207042, 266.522625215281, 
    265.109636815528, 263.698795848737, 264.018661381438, 267.888987960721, 
    269.85725104376, 267.763670176944, 272.912325403583, 277.725671690989, 
    276.323093039103, 275.868165753673, 275.018379214849, 271.790703278643, 
    266.535243162486, 266.851640834053, 267.202733242762, 266.580740612275, 
    267.418163055204, 267.42717884936, 267.066644188296, 265.42521342888, 
    263.530412460353, 261.812746028957, 263.770672200872, 265.382086596625, 
    269.769163845334, 278.244104645586, 278.438407098795, 276.254576897728, 
    271.513063075698, 266.541991288216, 267.810451906382, 269.526849536193, 
    277.311072376919, 278.506838397038, 273.677101091626, 273.618346761196, 
    274.189123698136, 273.541801582131, 273.92404873319, 269.177658637985, 
    269.559046544474, 269.236229292628, 266.432618388061, 266.988925803845,
  268.64664463561, 269.931869532856, 269.095990623954, 268.267385242788, 
    267.076902358644, 266.227488379651, 266.094553302645, 267.210515190345, 
    269.870956658623, 269.745144867384, 267.506083071085, 267.534453901947, 
    267.382168231436, 265.931338620877, 264.796243685001, 263.83443122458, 
    264.300465169131, 267.19589569899, 267.466042342294, 268.415795691906, 
    272.371193649247, 272.98654012294, 272.898180290187, 271.75710476706, 
    270.58455230615, 269.888371321752, 268.449823177902, 266.781553683493, 
    265.593397519815, 266.107891244973, 267.026932564668, 266.666697598469, 
    266.557743930421, 265.690208808873, 263.438306284307, 261.24489349069, 
    260.146795281053, 259.908266851662, 261.791129769684, 267.717194060832, 
    271.078503385658, 273.507731394335, 271.547572619622, 268.895111198654, 
    267.870979613137, 267.638691902977, 268.790649460239, 273.573808566374, 
    273.287605042857, 271.912556576676, 270.481056225488, 267.703172403279, 
    268.586806541241, 268.389767199008, 267.807166102986, 265.529507998352, 
    267.118678009107, 265.902744686906, 264.021039872398, 265.031356781405,
  266.10511833484, 268.447266645538, 266.373991657135, 265.656485179295, 
    264.287380079987, 262.724864820216, 262.052432863438, 262.344275185973, 
    265.111639446949, 266.894112115697, 266.006596831565, 265.704078416244, 
    265.619171303224, 264.597527182191, 263.895079064916, 265.281113704403, 
    266.200187898542, 265.791334661508, 267.518049190266, 268.354712744184, 
    269.39306474449, 269.17666632219, 268.323949824391, 267.068132667565, 
    266.427991963666, 266.044377988055, 265.39515063422, 264.845865171227, 
    263.949477061258, 263.638546788866, 264.263079541602, 264.67520696241, 
    264.778313575002, 265.280092747615, 265.980187956934, 263.483817657172, 
    261.740712026036, 262.984982138264, 265.670603833958, 269.642247193375, 
    270.105608763832, 271.285359785629, 269.641009392058, 268.324751684846, 
    269.444589372103, 268.465311485813, 265.567521098612, 266.49418077167, 
    271.758974562905, 268.712634164648, 267.065187673918, 265.525114582279, 
    264.089534631524, 263.553901226986, 263.517047592606, 264.157510740967, 
    264.861960750379, 263.745000881166, 262.647676783231, 263.722182217624,
  259.809810065712, 264.037459344726, 264.526528040227, 264.49899914488, 
    264.187827979446, 263.30622893671, 261.063429557127, 257.800952332329, 
    258.003864656365, 260.578788756912, 262.289654360775, 263.56053047567, 
    264.350789214343, 264.045546542876, 263.283866481706, 263.602409251688, 
    264.257932479585, 265.373678548646, 266.248656749213, 267.667747060762, 
    267.530853184801, 267.454120971129, 267.757483127891, 266.922207328254, 
    266.9954770393, 267.981245043277, 268.911163679811, 268.260114871866, 
    265.795163141774, 263.232507340461, 260.973413580579, 260.216403985697, 
    261.007916844899, 262.191528629422, 263.202393803319, 261.754111571471, 
    259.712469616388, 255.653170795971, 260.513996637104, 266.935389748067, 
    266.595716085197, 268.684685086621, 269.744693467218, 269.180599701435, 
    269.021222419404, 268.690244437718, 270.240364579737, 268.392016283826, 
    261.860139954913, 259.718690381775, 262.582136983651, 262.818005864978, 
    260.956252649801, 259.390182188021, 258.342120500698, 258.179641897157, 
    257.911318452926, 257.105204988699, 257.181802212139, 257.989094256381,
  256.664760674091, 258.407996996735, 259.922441799877, 260.992272800478, 
    261.705424623223, 261.556497463722, 260.574293873241, 259.209434520272, 
    257.239257424337, 255.226396697295, 256.091382527058, 258.465456203822, 
    259.858527461584, 260.358305405919, 261.004161613551, 260.566592171987, 
    260.09725583024, 261.586761322657, 263.535240569767, 264.781725374308, 
    265.722037660051, 266.284906962096, 267.444609989863, 267.713955819328, 
    267.055109916446, 266.591809309986, 267.53717033795, 267.406698317689, 
    266.114229671132, 265.643785540749, 264.535055187619, 262.898579024754, 
    261.680612745343, 260.644320597679, 260.308749645041, 260.234771895166, 
    260.00506169419, 258.646313326523, 258.899385173796, 257.197298166213, 
    257.623703934873, 260.36557403804, 262.083996928144, 262.328696735574, 
    262.637189551684, 262.965742021666, 264.171903080917, 265.4116084018, 
    265.148743788603, 264.633868726066, 264.104188188382, 263.433318940818, 
    263.453467666593, 263.43558008984, 263.053578819107, 262.432691346944, 
    259.929786024816, 256.634851943671, 255.892294524374, 256.433647065325,
  256.677043417057, 256.313419741492, 256.371824460991, 256.689583910584, 
    256.763575411078, 256.473207663975, 256.330434268072, 257.007993442625, 
    258.184843411858, 258.510249657914, 258.014421956989, 258.154795255556, 
    258.905664128509, 259.471192190968, 259.737125978164, 259.747371739319, 
    259.843193015503, 260.301242690838, 261.273702463806, 262.619344695381, 
    263.766760286263, 264.482087088844, 264.723524707801, 264.328278803139, 
    262.782373882066, 260.297730953697, 258.478136268103, 258.444474983549, 
    259.097650601143, 259.520917540652, 259.319903198358, 258.802088916101, 
    258.232915873536, 257.686648104091, 257.321054064477, 257.153566951847, 
    257.093553403777, 257.279947931876, 258.107384701055, 259.181903867724, 
    260.023568189036, 260.369201571021, 260.626898637575, 261.092111260785, 
    261.469773389069, 261.563004302892, 261.611231310164, 261.604227166534, 
    261.640607651827, 261.408663385095, 261.671543492992, 262.405162164258, 
    262.58154860468, 262.15756646934, 261.544558557617, 260.873111796835, 
    259.044886612474, 256.939986465135, 256.696753150985, 257.089682876888,
  257.147443096682, 255.835142945702, 254.746644365301, 254.1439442499, 
    253.903051727381, 254.252603656756, 255.106557290287, 256.049706347632, 
    256.665728914819, 257.017362179121, 257.285582241399, 257.500262919745, 
    257.570304892568, 257.47094311364, 257.407048838742, 257.447892714299, 
    257.52778293671, 257.696427168157, 257.975666407439, 258.236962217125, 
    258.538250047131, 258.85136785033, 259.025625017266, 259.124140338632, 
    259.08049467286, 258.937685599719, 258.948230347948, 259.013055762436, 
    258.918515114103, 258.705714128787, 258.412470213114, 257.982753941081, 
    257.528373220657, 257.140616573296, 256.86652826629, 256.767409067637, 
    256.840713380083, 257.036939350675, 257.299657492014, 257.746742063002, 
    258.144645590279, 258.281718336261, 258.294516219256, 258.349422941579, 
    258.318447847937, 258.256851362695, 258.222776519733, 258.236138297019, 
    258.290259213234, 258.314076053897, 258.427098627269, 258.463707486505, 
    258.406945758561, 258.417795854832, 258.407746575146, 258.299256894466, 
    258.057187101006, 258.031450816793, 258.225101694805, 257.990971982442 ;

 u =
  8.84831659633795, 8.77622627592505, 8.74661515523524, 8.80012838018033, 
    8.95262292826209, 9.21712610781407, 9.5825750551377, 10.0129219981738, 
    10.459243214595, 10.8692440542647, 11.2035086077027, 11.4455857127763, 
    11.6015855607979, 11.6844679703426, 11.7032665689987, 11.654826203879, 
    11.5624237917244, 11.4138648685502, 11.2383118647152, 10.9907716743336, 
    10.6444657717831, 10.2213426206817, 9.7420337981308, 9.22046836987497, 
    8.6827193948523, 8.17903579157798, 7.76089711905612, 7.4388415264334, 
    7.23130367585518, 7.16233515453806, 7.21753680677805, 7.37024045846886, 
    7.62301900269402, 7.97509501446704, 8.38942311997003, 8.81800127834139, 
    9.21428152605042, 9.54459333804197, 9.78653192384891, 9.91484294820113, 
    9.9299406320172, 9.87280083630531, 9.79591089095981, 9.69372303484705, 
    9.57507553049623, 9.52367876388992, 9.56057205457846, 9.61384531227116, 
    9.63828651857039, 9.63606554996548, 9.62154869737901, 9.5930403592359, 
    9.53623694885524, 9.45757788279343, 9.36845445788878, 9.27609308816585, 
    9.18854300161254, 9.10486722458318, 9.01767360778439, 8.93142588589542,
  7.41851788587563, 7.33976839931418, 7.30184151091704, 7.34562579349439, 
    7.52701623985026, 7.81821248906549, 8.16825875912297, 8.59770185939013, 
    9.11489863248394, 9.65858973306529, 10.1174880572904, 10.4123166351743, 
    10.5134710329851, 10.4779337208722, 10.4031188866668, 10.3590549539869, 
    10.301251777803, 10.1996089124456, 10.0817427812504, 9.98102192895391, 
    9.8085530773114, 9.50966685528361, 9.07508211352004, 8.57582507714715, 
    8.11317189781143, 7.69471485007376, 7.32822179652016, 7.07110752340417, 
    6.8764127640774, 6.71982672399787, 6.69825249510421, 6.80914660337965, 
    6.92013427354873, 7.03757269617282, 7.21693312604188, 7.4343272644059, 
    7.68489175940596, 7.9731523530246, 8.23331311193606, 8.40033338880308, 
    8.47550782398553, 8.48279871084076, 8.44391736212012, 8.37883319534577, 
    8.27308712892157, 8.17525310490646, 8.18563590941968, 8.30471701529392, 
    8.46384054167488, 8.58124186888431, 8.62010271106943, 8.59062160441584, 
    8.50415071294039, 8.36640714923242, 8.22069707587903, 8.10415583431617, 
    7.96909857706392, 7.83427992366108, 7.70054123324487, 7.54616427567243,
  6.6417776743045, 6.52225186586992, 6.40903964407888, 6.26073542524193, 
    6.2061873025234, 6.30108474105196, 6.54610907480549, 7.02921396545942, 
    7.66517780759436, 8.34612435708113, 8.95724037834359, 9.42621031869329, 
    9.63382744388348, 9.53788266108842, 9.32124533978495, 9.11138420040117, 
    8.9537409309506, 8.90965628922274, 8.93596834050448, 8.90647179528525, 
    8.87658619710778, 8.86658110916319, 8.70246228242438, 8.28033018690646, 
    7.75035715841419, 7.35734725643206, 7.09043338447723, 6.88030061380816, 
    6.83371134398398, 6.81323591091645, 6.75066388430248, 6.76437799872472, 
    6.84302566950615, 6.83127053980793, 6.76174225548834, 6.74064445495803, 
    6.86264832718704, 7.02536549154538, 7.13207861322974, 7.20537160366533, 
    7.28456843074526, 7.32806624305605, 7.32165394088214, 7.3083492954602, 
    7.27350396960997, 7.24059370081894, 7.2400226650799, 7.2936383570425, 
    7.45189388253564, 7.70899806977759, 7.9088165031204, 8.01094218126012, 
    7.91480166636121, 7.76836663355051, 7.54294460426676, 7.37275748085655, 
    7.19888818830869, 7.03672802610905, 6.93194990857183, 6.80290772924849,
  6.11609077542862, 5.98478699260759, 5.77319261768944, 5.4958275688978, 
    5.17356707333524, 4.93040880970401, 4.89674498670565, 5.14042901319283, 
    5.61937781997683, 6.22424057537666, 6.78200925843609, 7.2999717850563, 
    7.77127854441901, 7.826268556125, 7.52231118070854, 7.01565482029581, 
    6.60488004811595, 6.51658747297679, 6.83189007113144, 7.10287066517934, 
    7.32680446547454, 7.4346020441929, 7.37351728688514, 7.08977322150249, 
    6.72009649909884, 6.46162352858061, 6.33284948664549, 6.2128768220587, 
    6.21679274307074, 6.53058302211555, 6.75946117539282, 6.7626769859991, 
    6.71864633324772, 6.6328000940924, 6.31186087835347, 6.0658107865715, 
    6.05274467458172, 5.98166068403762, 5.88529665499231, 5.93439392506334, 
    6.08337366594515, 6.17305889963997, 6.1587104729561, 6.08596753236175, 
    6.00733395025749, 6.03540533919011, 6.16491604469559, 6.2460440632147, 
    6.32719557855312, 6.57853346063741, 6.69935380248358, 6.84504346148486, 
    6.80329051499779, 6.73929314148874, 6.60638469744009, 6.2093953145007, 
    5.9349471216551, 5.85497482580137, 5.91818659017714, 6.07762523981078,
  6.02738107894249, 6.0063223288964, 5.86376837050585, 5.62126980195601, 
    5.24786115513758, 4.84174784973322, 4.5885910170664, 4.43379726907497, 
    4.41741919779126, 4.65492622276087, 4.98994743907692, 5.42976623548951, 
    6.08552340935682, 6.30286485368531, 5.76165149865893, 5.08190071407795, 
    4.64140371593572, 4.44779102975643, 4.78143819964455, 5.36946772693231, 
    5.94032733756258, 6.20398615248231, 6.19878007880514, 6.00022691138727, 
    5.80243353672429, 5.62487483766425, 5.57863600947694, 5.65352915412819, 
    5.7531025660097, 6.10603589359048, 6.53415409539369, 6.94852868335438, 
    7.05061037026487, 6.85575166515881, 6.33301482051832, 5.87098865502915, 
    5.59833854502578, 5.38992417252944, 5.36948572309982, 5.52838556506477, 
    5.64758935705904, 5.6419851277298, 5.52429388662665, 5.40597016628207, 
    5.42174398359073, 5.55901307695726, 5.7729678818253, 5.89364352339725, 
    5.95982654477895, 6.09529188662914, 6.01977764820495, 6.09402461151203, 
    6.11171437210731, 5.84644108465078, 5.63567756707623, 5.23024983229665, 
    5.05477468597214, 5.21811647533537, 5.49077824225529, 5.82548827250383,
  8.33557483594457, 8.56083888244734, 8.41462814089551, 8.11598750163753, 
    7.8136484493305, 7.46598602661247, 7.08176323204516, 6.6760061737491, 
    6.30696956162869, 6.03223157066214, 5.96062452337106, 6.13362250636991, 
    6.71648464201056, 7.38315010165398, 7.0403017577819, 6.00859721176617, 
    5.22061946534933, 4.85119795839613, 5.15921809007909, 5.98426580320452, 
    6.81991174150477, 7.55572793437009, 7.88270146234284, 7.79273577836181, 
    7.61074844676592, 7.54048511156064, 7.47790355200899, 7.2908749414505, 
    7.36195703644192, 7.57347812406708, 8.04919767174314, 8.77584986571494, 
    9.10940705450612, 8.77935648428277, 8.27605358129327, 7.81352600608127, 
    7.44173749399338, 7.21059726324642, 7.24747835508666, 7.49145023696662, 
    7.7017161396873, 7.72667345719696, 7.52805532360484, 7.25544002043655, 
    7.11528937918895, 7.18426239562787, 7.47328339429874, 7.84814070645326, 
    8.15432507150709, 8.08180698697888, 7.76558705880398, 7.72737298005465, 
    8.03357698127478, 8.05709764526883, 7.34370771752718, 6.67289511026459, 
    6.52232950259517, 6.72224174247565, 7.13390804867113, 7.75575093943376,
  11.5466375923218, 12.3018221026398, 12.4306737627108, 12.1275663804487, 
    11.670562447397, 11.3244628193235, 11.0718360975898, 10.6469515843619, 
    10.1005502248348, 9.48405084885744, 9.04770321589169, 8.83350982189489, 
    9.03907604971332, 9.69956282025099, 10.0740668630852, 9.58957529483345, 
    8.40294264264672, 7.48275095127379, 7.37207230714482, 7.9491047513525, 
    8.92082217562885, 10.2497140087866, 11.3108154083716, 11.6099448934052, 
    11.4464791251677, 11.2242460242144, 11.1189904483574, 11.0560957712099, 
    11.1767452616434, 11.0946455452588, 11.3257903508424, 11.7387365436505, 
    11.9355112808269, 11.5994222225811, 11.3419979408328, 11.3086118984369, 
    11.2792944953394, 10.9246458942784, 10.5778340938933, 10.5513934982137, 
    10.8484289495421, 11.2103436468884, 11.2621949576415, 10.9476053979408, 
    10.4323616232395, 10.0541654751919, 10.0773693157477, 10.4885543030261, 
    11.1764138144126, 11.5073555167323, 11.2491454093299, 10.8513784990105, 
    10.8853022360541, 11.5241330720147, 11.6620143265983, 11.0605973035151, 
    10.2704305265525, 9.75236076910352, 9.82742219859279, 10.5512089195994,
  15.3574574582778, 16.6398923240828, 17.2260256071526, 16.9911872135697, 
    16.4004731323613, 15.9033702632637, 15.8788160446956, 15.7656962457875, 
    15.2662257177535, 14.6186486763117, 14.0345869779463, 13.5817647295541, 
    13.3632809073538, 13.5227003145416, 13.9862384185853, 14.4227423736101, 
    13.9219541511494, 12.8865042957873, 12.0126185482949, 11.9311129241594, 
    12.6281890516461, 13.8721822358735, 15.4818001321554, 16.5875668626739, 
    16.5994488704941, 15.8104550556359, 15.5348750963164, 15.8217154885886, 
    16.3511625004747, 16.7109359518018, 16.7782697939189, 16.2131739368829, 
    15.6177557760597, 15.1430600057813, 15.0612662140896, 15.5322828436049, 
    16.1288068598432, 16.1709327469549, 15.6401266306801, 15.0258215823439, 
    14.9123473786011, 15.3792418189935, 16.0170017961495, 16.1002146342957, 
    15.4171692551582, 14.5968480547813, 14.0942644500322, 14.0884213701126, 
    14.7181814418206, 15.4728014284013, 15.7893019058318, 15.3476244340211, 
    14.8518701412115, 15.2269625464474, 16.3599847130479, 17.0488001321742, 
    16.4223214903326, 15.204522335886, 14.3934849670364, 14.4954352111027,
  21.6514094444324, 23.0644759342539, 23.8844535510542, 23.686545169203, 
    23.0887551341184, 22.3980522853207, 22.4782868140009, 22.6481518208861, 
    22.3800764223976, 21.9360757992244, 21.356329666577, 20.9251768272876, 
    20.5981197300107, 20.4727962451674, 20.6980535532501, 21.2210515820564, 
    21.5419638188488, 21.0592331581921, 20.0702173785897, 19.4607979863878, 
    19.6245098527143, 20.4530481006847, 21.8830835899643, 23.4103526358303, 
    23.4971136333398, 22.3798197705659, 21.8778387843207, 21.9724278908956, 
    22.744029486472, 23.8248207003426, 24.2807126543979, 23.3928099353276, 
    22.1554888465306, 21.284702955788, 21.015839068588, 21.4821639367516, 
    22.3956081421604, 23.0974637369392, 22.8867387761916, 22.0324297832186, 
    21.5429914693546, 21.7749218638264, 22.648558877424, 23.3240753461508, 
    22.8519695509209, 21.8627653499069, 20.9400748585201, 20.4982334325534, 
    20.8634854871055, 21.5801196954837, 22.1223869536947, 21.8157029488182, 
    21.2549938558219, 21.2369478423559, 22.1767641544509, 23.7824520913396, 
    24.2987145531409, 23.2548722303318, 21.8382447789408, 21.2345718088161,
  28.1897981552393, 29.3395789055118, 30.0403330722387, 29.8371602730645, 
    29.3120183364763, 28.6363599741152, 28.7360195407238, 28.9977033123651, 
    28.878378256487, 28.5932086325274, 28.0793178737632, 27.7747919601972, 
    27.6527177664314, 27.5132667092197, 27.6736592553265, 28.0824477781331, 
    28.5356909174254, 28.2395461135867, 27.6974614320145, 27.1756118381942, 
    27.0409908049692, 27.6012917689387, 28.6530357394367, 29.8875140923651, 
    29.571296562353, 28.6522953018546, 28.0415306903548, 27.8563434785936, 
    28.5468773652676, 29.6790196795643, 30.4011086250659, 29.8997972898179, 
    28.808515120214, 27.8260956249267, 27.39638067723, 27.5738092873368, 
    28.4729684319498, 29.3527124357866, 29.3423523837774, 28.6267317114587, 
    28.1104120821707, 28.2196837611456, 28.987739894359, 29.8128998236572, 
    29.6470726222832, 28.8648377443508, 27.9058097722204, 27.3132565661787, 
    27.3663937255597, 27.917235516735, 28.2924293625368, 27.9128631488713, 
    27.5061232549064, 27.3629405220339, 28.0350474028911, 29.6459742887688, 
    30.6644560573057, 29.9936208837417, 28.7560659935385, 27.9982550836926,
  31.8092314843884, 32.5713770567093, 32.8374780227591, 32.5630414286106, 
    32.1761050188828, 31.7854872469206, 31.8731666856915, 32.1609052261193, 
    32.0710120955715, 31.7440748012753, 31.3009787250072, 31.1912808862355, 
    31.3103997850636, 31.4741082498317, 31.6682793697026, 31.8847932342967, 
    31.8091988646208, 31.6029672208559, 31.3940315006411, 31.3292515777208, 
    31.4236949204934, 31.7358298036263, 32.4374229458359, 32.9807125005779, 
    32.26089210418, 31.8142399387956, 31.1861426700842, 31.0354132952221, 
    31.6657194985082, 32.3091259700978, 32.7083155196686, 32.5852611627549, 
    32.0623761841374, 31.3024499114265, 31.0699538408471, 31.0502163200065, 
    31.7853592435012, 32.4631779672644, 32.3470359783157, 31.8946358794564, 
    31.5092621485825, 31.6495818585534, 32.3316003567482, 32.7159946602973, 
    32.6744862873711, 32.2296888605118, 31.6078398889363, 31.265168383223, 
    31.1517084849693, 31.4693109123177, 31.5365705371619, 31.0288996724743, 
    30.8474021767821, 30.7008514661052, 31.4002184947809, 32.7113372826107, 
    33.266378020445, 32.746680347478, 32.0498437619477, 31.5235128650046,
  33.6267949359107, 34.0112638630451, 33.8783003367787, 33.5275021046701, 
    33.1282944553235, 33.1837354128381, 33.2967068591435, 33.5808870421096, 
    33.3568867166351, 33.0803967956042, 32.731629968382, 32.8631877414055, 
    33.2269751084501, 33.5738295990671, 33.7874774965444, 33.7548863216078, 
    33.1204603592971, 33.0909211319376, 32.9996381955245, 33.1758257490105, 
    33.8766428113984, 34.0334880068062, 34.2230333636204, 34.0389767464932, 
    33.3636342782538, 33.3173568080922, 32.9132712382894, 32.6938532486338, 
    33.2710404976224, 33.6383017614229, 33.5664100307764, 33.4737098944891, 
    33.4044683504962, 32.9308933349482, 32.9336221964045, 33.0172218736014, 
    33.4337488051597, 33.7873068925791, 33.6319252193878, 33.4031624023501, 
    33.2419090108928, 33.3290752696271, 33.7869535865656, 33.8627072573741, 
    33.7817392267511, 33.5162885516177, 33.2237080484535, 33.2001304337167, 
    33.2058454222246, 33.2562483841813, 33.0897027292493, 32.648833899006, 
    32.5900852851854, 32.599945915978, 33.3413478493757, 34.2317142719232, 
    34.2236759933289, 33.7418504201932, 33.4893551951521, 33.2875989895895,
  34.2236926359789, 34.3849417085985, 34.1775967818494, 33.8435952000352, 
    33.3738800766683, 33.6995742929869, 33.8664716827201, 34.05145962186, 
    33.5663807742254, 33.5817822665379, 33.5826962815286, 33.8541155209052, 
    34.26487896661, 34.5148477831586, 34.6029146061426, 34.349526891535, 
    34.0777267619154, 34.0974587745031, 33.8156382645663, 33.8537502799632, 
    34.9453795885494, 35.2075774459463, 34.8156383133951, 34.2124862902553, 
    33.9863778418747, 34.1270768354225, 33.9434473463332, 33.5629773746125, 
    33.8731164791382, 34.2020192391302, 34.0113603756115, 33.8184099737466, 
    33.8903051442189, 33.6881799391523, 33.7381510617831, 33.9770410291335, 
    34.0919697636248, 34.1667637908838, 34.1320200597505, 34.0593775077805, 
    33.9523053643997, 33.9721040657681, 34.2698601018555, 34.3359080686867, 
    34.1743451908274, 34.0642317358082, 33.9213284744293, 33.9683083191815, 
    34.0686709859075, 33.9439616783057, 33.7742873230198, 33.6312098900539, 
    33.6934203280666, 33.7452111396785, 34.213210177704, 34.6819672863002, 
    34.6705788388776, 34.2626132631793, 34.2402769844237, 34.1791658658745,
  35.2845048667323, 35.3034195173057, 35.2042604259847, 34.9057834724433, 
    34.6404615318639, 34.9609654073825, 35.1640536163188, 35.0829948880274, 
    34.766944714657, 34.8420196847613, 35.085721903499, 35.3425557776509, 
    35.6111175488557, 35.7558326818756, 35.7319948436359, 35.4926448155487, 
    35.8667393251092, 35.89046228173, 35.4842021341652, 35.3745610016953, 
    36.040706858554, 36.367473979818, 35.9295587752252, 35.3702989461194, 
    35.5032141922567, 35.6558188875243, 35.455702819951, 35.2792329942655, 
    35.2137013676491, 35.3559500852002, 35.2284253852018, 35.0186919182564, 
    35.0501530775627, 35.0589375148761, 35.0907381254319, 35.2720086119374, 
    35.3249792533434, 35.3253753408289, 35.2920568783165, 35.2940470742256, 
    35.1526650557673, 35.2550153734764, 35.5395463558567, 35.4767028796344, 
    35.2766056653561, 35.3384317860941, 35.3280007934739, 35.3609522960675, 
    35.4331329852142, 35.2624068928824, 35.0348129240621, 35.2907886471369, 
    35.5596117247212, 35.4755683880805, 35.5609940154014, 35.8016216668784, 
    36.0255548326946, 35.7484440591318, 35.6650795833275, 35.5767490536499,
  36.1982738789347, 36.2974746232973, 36.1096130444223, 35.7517822694473, 
    35.8657299074653, 36.0616627607662, 36.2320704653926, 36.1156987664279, 
    36.0340148061015, 35.7518067752093, 36.0781530900417, 36.3569084693159, 
    36.5342868344121, 36.6702502164743, 36.6581299232838, 36.5766437213558, 
    36.9619124790017, 36.9072649921227, 36.7772629902165, 36.7786200785558, 
    36.8316328452103, 36.8925448313665, 36.7915603325391, 36.4530976494515, 
    36.63385149624, 36.7563772835574, 36.5718834034647, 36.6865366259648, 
    36.3552302431662, 36.2972066418341, 36.2364837953304, 35.9857874997705, 
    35.9676320087678, 36.0802538895736, 36.0988926623637, 36.1596808711984, 
    36.2538230391695, 36.3186197517451, 36.1909789436521, 36.1176574730525, 
    36.126764425171, 36.3301987767204, 36.4603215590385, 36.2394533360156, 
    36.1255956378148, 36.3365297346651, 36.3879439774302, 36.4727130404561, 
    36.6401993985166, 36.4577131639115, 36.0684594992161, 36.4998499959132, 
    36.8707310705036, 36.7876313612608, 36.7112700374929, 36.8091632973928, 
    37.092731879094, 37.1431654221936, 36.7198351705216, 36.1256421368876,
  35.3834917807553, 35.5700718231753, 34.9997350525198, 34.5865176190962, 
    34.9389318611161, 34.9772592941381, 35.0621487222951, 35.3097957829554, 
    35.2562736941587, 34.9158467326788, 35.1401861419746, 35.2839549544325, 
    35.450872484469, 35.6013323062466, 35.60954033494, 35.6581624588669, 
    35.7884909094305, 35.6937012571905, 35.8391742965638, 35.8648132378351, 
    35.7911941624129, 35.6734528973446, 35.656451451917, 35.3636473241469, 
    35.4674586071339, 35.6474706340087, 35.6982401812082, 35.8326157495241, 
    35.4902106942566, 35.3587905548588, 35.2761040579322, 35.0756279758552, 
    34.9810373012928, 35.0131310900506, 35.0173997831407, 34.9818468870805, 
    35.0784546028798, 35.2107284814367, 35.0806122973084, 34.947659467153, 
    34.9966262071863, 35.0950998942656, 35.1150491357678, 34.9999576186552, 
    35.1385967586606, 35.4158081331937, 35.435498657977, 35.5161241937764, 
    35.644211121025, 35.57461165238, 35.3732918884888, 35.6780323213824, 
    35.8674080497857, 35.867053599375, 35.8078692620932, 35.8226213450369, 
    36.0142018575971, 36.3824330858208, 35.786387332036, 34.4466579310155,
  34.1677216465415, 33.9988180123636, 33.2135396470328, 32.8313098166578, 
    33.1265875792267, 33.2193230664358, 33.4895736223087, 33.8757841360492, 
    33.7804784421319, 33.639396622477, 33.5919301028024, 33.6077847223436, 
    33.7167521663665, 33.7655585362755, 33.7913753507142, 34.0337274883858, 
    34.2198466153318, 34.1414492189955, 34.2063674662171, 34.1683974049557, 
    34.2411257781512, 34.171074919882, 33.9322800334243, 33.5246866722691, 
    33.5894780312908, 33.8849137626894, 34.1983967658282, 34.4027507541783, 
    34.3442165428492, 34.2731131960484, 33.863088400307, 33.5696675427468, 
    33.2960303585125, 33.2468904921817, 33.3582648807082, 33.3450818483796, 
    33.4432029790664, 33.5610138647179, 33.3973143480849, 33.2043756147056, 
    33.0830252523634, 33.0444473562107, 33.1194472806054, 33.3459586944306, 
    33.7993231411846, 33.9674453283242, 33.8615914072192, 33.9078779214983, 
    33.9175136862177, 34.0206670082209, 34.1705148117735, 34.3166740479113, 
    34.2630890962135, 34.2662235764907, 34.2964729144674, 34.3865307710428, 
    34.4109850587785, 34.6804503427872, 34.2818296054642, 33.1590574380577,
  33.1974265868594, 32.7737689693677, 32.0993398945631, 31.7152846684573, 
    31.7326598529381, 31.9922063263929, 32.6839465975735, 33.0959827197054, 
    32.7060340254165, 32.361390702786, 32.0783817528556, 32.2278808995544, 
    32.4074429364746, 32.4043155575708, 32.4777304867146, 32.9073011450353, 
    33.3027686040254, 33.2003510992877, 33.0457395107653, 32.9051628525701, 
    33.1322819530362, 33.2165551429298, 32.7771065613602, 32.2712139680978, 
    32.3341580795544, 32.702604191233, 33.1554199554216, 33.4882543505526, 
    33.6558494776378, 33.7361988245168, 33.0571790686068, 32.4777247296754, 
    31.8520144006848, 31.79136075152, 32.1397072209842, 32.2414921179924, 
    32.4692603930043, 32.6206804733098, 32.3194609251099, 31.9116869463799, 
    31.513358702342, 31.3774136804403, 31.5660315709887, 32.1202361325064, 
    32.80442042353, 32.9810984561893, 32.7846994120384, 32.8256487794523, 
    32.9384960950636, 33.0782150808697, 33.2346622252642, 33.3157861423932, 
    33.2478250396185, 33.1826424975674, 33.4150491540531, 33.7070170867117, 
    33.4571863144912, 33.3894231363795, 32.9802334318864, 32.7175757093737,
  31.0411117536373, 30.8378275778209, 30.2808626515001, 29.7630899299429, 
    29.4040583529131, 29.668497763861, 30.5382343241665, 31.2598459542233, 
    30.7460591392722, 29.9845781680395, 29.3429121032733, 29.2625877369055, 
    29.7828701464415, 30.2904711632069, 30.7169393925606, 31.1900735966039, 
    31.3817195245729, 31.0876499392377, 30.8227450859564, 30.645979734282, 
    31.0862659742291, 31.1841600678016, 30.6680386716722, 30.1983328945517, 
    30.1731784960836, 30.5555806262294, 30.9814378856777, 31.3115445995481, 
    31.5405402493566, 31.7567208350899, 31.278447230686, 30.5193413880999, 
    29.6315338096036, 29.3662639048518, 29.6514636092302, 29.8804742645865, 
    30.4592947168679, 30.9021442765059, 30.522555086782, 29.7642888815307, 
    29.0190902154435, 28.6561147959917, 28.9224654663224, 29.6814132166597, 
    30.5079826849944, 31.0079888437273, 31.0180774667731, 31.1138014126999, 
    31.1793561344535, 31.1502724633099, 31.1612494140025, 31.091934270867, 
    31.0710089607806, 31.0406320020252, 31.4664908522498, 31.9226235898442, 
    31.4843468167788, 31.1540861945744, 30.6073932345272, 30.6425748062822,
  28.02966093333, 28.1089202265836, 27.4622796228105, 26.8054703572506, 
    26.1860335804745, 26.3623796840679, 27.2363609219138, 28.3195034848984, 
    27.9923328266223, 26.7298334153774, 25.7179909661894, 25.2198828269589, 
    25.9802469323766, 27.4581430203799, 28.6634753941352, 28.8940162728631, 
    28.3798926383294, 27.6722971826112, 27.3602334170016, 27.4465487421143, 
    28.1651325713249, 28.1339134319765, 27.57687056942, 27.0393511088554, 
    26.6874602106361, 27.0337111637052, 27.5207825161909, 27.9423769056367, 
    28.2581220157111, 28.5466610999547, 28.4142724797775, 27.5228274820517, 
    26.5579882246902, 26.0915354586018, 26.1935940091181, 26.6671076845978, 
    27.7950894129216, 28.6587763963905, 28.114491543613, 26.7832312331086, 
    25.6271530484887, 25.0680712257604, 25.3661999378921, 26.2806002673194, 
    27.3414067912104, 28.267039971939, 28.5579234976104, 28.5100510499451, 
    28.2675696459073, 28.0062086695242, 27.8829515411382, 27.700245376926, 
    27.6578478760107, 27.7456262949318, 28.1916623680448, 28.6899728458325, 
    28.4605987994562, 27.9125979465793, 27.5277733200279, 27.5061283476351,
  23.5056952050142, 23.4980747625455, 22.6976571955028, 22.0981355015966, 
    21.7806177646193, 22.0592710770046, 23.0324867167427, 24.2352696172068, 
    23.8376971318488, 22.0916215113299, 20.8528859734037, 20.4476360405757, 
    21.4721241858212, 23.6284282318454, 25.2523650043847, 25.0592354537136, 
    23.8751858340852, 22.8256401721568, 22.5210165411074, 22.898902248979, 
    23.6853584021355, 23.5945538372048, 22.7817385949576, 21.9954735725789, 
    21.4779680695679, 21.7584318824462, 22.6078101140946, 23.3298850553965, 
    23.6844736788514, 23.886041909944, 23.6880195706078, 22.6904126764451, 
    21.7979908608828, 21.5852586741568, 21.9090691223988, 22.7783906476074, 
    24.3625589459942, 25.1365759706916, 24.0990287993872, 22.2151774004208, 
    20.8493036623964, 20.3299942467077, 20.7601612931363, 21.8354527895484, 
    23.1870615492554, 24.2714914099397, 24.4366125180218, 23.9435470140989, 
    23.3654204605049, 22.9700695188054, 22.7256010996166, 22.5545860639428, 
    22.5102741140821, 22.6124413909443, 23.1405631601222, 23.8167259720824, 
    24.051397166367, 23.5332550703708, 23.2551917620576, 23.1616470022807,
  16.1547104718441, 15.9844354033517, 15.6676807141758, 15.6591089684647, 
    15.9452177218734, 16.4605431237254, 17.5379768724423, 18.3173447921958, 
    17.329445252591, 15.5366998766212, 14.6146525293635, 14.8361463727624, 
    16.2421069965156, 18.281574704653, 19.329664042792, 18.6972238958335, 
    17.3050548754556, 16.2579910722014, 16.0185698529098, 16.3092249270258, 
    16.7405027853222, 16.4600294646309, 15.4213703451974, 14.774070288274, 
    14.593041271285, 15.0319050153152, 16.179475171549, 17.0225929587707, 
    17.2584784581842, 17.0905445774097, 16.4843526474918, 15.6622951965904, 
    15.263935488247, 15.6107824855613, 16.4791677755736, 17.8620400750027, 
    19.2090209044821, 18.9576134314414, 17.3687453167933, 15.4857185984822, 
    14.3492313884966, 14.1199619936779, 14.7107173206075, 15.8628357802034, 
    17.3036262528115, 17.9972799686336, 17.5153150392725, 16.6128635918443, 
    15.7828721021995, 15.3988329635309, 15.2836060043545, 15.2903740720734, 
    15.4966026630705, 15.6725566724652, 16.3359954223969, 17.335898483433, 
    17.8318688361664, 17.421258907835, 16.8450980217708, 16.2765821484831,
  10.8370058072793, 11.2648976455761, 11.8081121398667, 12.2583973384297, 
    12.9370004790581, 13.7650099169357, 14.2583666952243, 13.929392246155, 
    12.7274647105736, 11.6330385029219, 11.4621183896694, 12.2790667802547, 
    13.6373878633578, 14.7539727656325, 14.8003271991071, 13.8556922072581, 
    12.6520642546438, 11.8314915608225, 11.6156943808725, 11.5434703517262, 
    11.394181669083, 11.0489939369767, 10.5226603423328, 10.568248664747, 
    10.9638016952023, 11.6355502032059, 12.5233571497462, 13.0107400237608, 
    12.9214997895959, 12.4069020568104, 11.8029408361136, 11.4759743838532, 
    11.7231660685737, 12.6382434626943, 13.9225770759238, 15.063544570101, 
    15.164982151236, 13.9024587657289, 12.3230763728284, 11.0319592213234, 
    10.3637340758336, 10.4866089923227, 11.300944338875, 12.488708209581, 
    13.3625624659633, 13.0626504738698, 11.9061998528315, 11.066154759391, 
    10.6566895653113, 10.5608726850816, 10.6328287739065, 10.8904365465623, 
    11.3001790931402, 11.7301943802922, 12.5297454122185, 13.4469708254784, 
    13.7171556977593, 13.1130113372436, 12.0892517302442, 11.1340797276061,
  8.01528837168651, 9.03614714566218, 9.83323220939153, 10.2744665677768, 
    10.8918311319652, 11.4206101482288, 11.0357766106772, 10.1979694320185, 
    9.62362055614199, 9.43262077388851, 9.76748064088863, 10.5038839268711, 
    11.169158754791, 11.2464227650512, 10.6501608601921, 9.68633304742709, 
    8.78065563075436, 8.19468351921672, 7.92403338124097, 7.72742994508681, 
    7.51267249156515, 7.65994494113466, 8.1019320843, 8.62325438635224, 
    9.13484191065569, 9.63010678649897, 9.97089514376555, 9.97025714307398, 
    9.62901294549441, 9.1953426728294, 8.92210326990375, 9.0256644330771, 
    9.72070534910624, 10.7293467416169, 11.4661290115854, 11.4774970762513, 
    10.6504890263171, 9.53007344623837, 8.5250167641046, 7.97919450779945, 
    7.86293217162297, 8.40503890658831, 9.36465078003638, 9.95286690059369, 
    9.68490994534069, 8.75334262062698, 7.74595198521191, 7.56173446828114, 
    8.08907561436346, 8.14926875378229, 8.05266077441815, 8.3973444890016, 
    9.00387309140344, 9.66208862635314, 10.2614592483401, 10.5159296664631, 
    10.3661992002326, 9.73956907054264, 8.76442736815115, 8.0164393672583,
  6.48893915911876, 7.23271694603013, 7.8783624870069, 8.30103183126553, 
    8.5413642460096, 8.47952142767789, 8.05859852314219, 7.60119290336917, 
    7.39734269335977, 7.45043715446948, 7.81145006108103, 8.09125254258665, 
    8.05983316926361, 7.66915128668036, 6.94312305820976, 6.18757797800528, 
    5.59673477715203, 5.2748126455583, 5.16331726971304, 5.21604394113668, 
    5.5095064747972, 6.11100622264364, 6.78718031030263, 7.20608673025216, 
    7.44770686747308, 7.61132356310599, 7.57114847950559, 7.29906362239168, 
    6.97332803656513, 6.75078742895759, 6.75070181478664, 7.06859883121854, 
    7.5750443235616, 7.95797664233915, 7.99645407957411, 7.53199835926115, 
    6.73735221094644, 6.24271573259261, 5.81936218495499, 5.80052527683351, 
    6.22459127879678, 6.95746535051696, 7.37336806563727, 7.12458657801886, 
    6.56799696696969, 6.06842629103158, 5.78031345587535, 5.87791330588696, 
    6.31559882756915, 6.36940730865187, 6.3845271296137, 6.66943254887421, 
    7.12993850216393, 7.51354101462789, 7.72058165227487, 7.70150222051049, 
    7.44933792232809, 6.98122124615348, 6.57060264585559, 6.25283191505192,
  6.06412588931154, 6.37685761985219, 6.76999105146123, 7.09684945365773, 
    7.21153084106374, 7.00839556891734, 6.72216880824425, 6.55943051244439, 
    6.49470134002449, 6.44065609584705, 6.45340967261322, 6.41644032863985, 
    6.24088320167146, 5.89380858291501, 5.38085933217876, 4.90809860015873, 
    4.59064719360895, 4.4982158703362, 4.68473507874549, 5.05018556290527, 
    5.62333552433451, 6.14297463262393, 6.47989049741614, 6.69312587737733, 
    6.76001787634272, 6.65376043737509, 6.41081379086872, 6.12086003147494, 
    5.87099724073269, 5.73666892454706, 5.78219410402599, 5.91114579613387, 
    5.92901477353298, 5.93768239657262, 5.95740944976816, 5.72750302086512, 
    5.31902563304546, 5.22285051121286, 5.27824841026882, 5.61356601953668, 
    6.17212396602728, 6.55801236536102, 6.57611306871454, 6.46049841591696, 
    6.29437704417776, 6.0967828498065, 5.93169605393963, 5.73270683570307, 
    5.64264416969169, 5.79528492667736, 5.97343230176955, 6.10089080160415, 
    6.16535557013493, 6.28078868380435, 6.41781904753178, 6.36119661409232, 
    6.13426355294487, 5.85523978329909, 5.83555125438706, 5.84909004062533,
  6.70466711892107, 6.82800627854234, 6.97133691534146, 7.11500574260973, 
    7.17823201580038, 7.12490802901039, 7.02607281464452, 6.92580100283945, 
    6.83015890757431, 6.71094780905864, 6.58220280201778, 6.46690578702724, 
    6.32116620991163, 6.09938557103679, 5.86705339058085, 5.73564925932925, 
    5.7453037865107, 5.85669070045046, 6.18211581490371, 6.62476577667844, 
    7.03546446532579, 7.31312372841733, 7.48331570327812, 7.55817835269872, 
    7.49884107732688, 7.2867156227945, 6.99603833003133, 6.73536635805154, 
    6.50828546331169, 6.28374550495291, 6.08361709533114, 5.96762693118664, 
    5.94904306674981, 6.00222617697334, 6.06476806515897, 6.14969221058948, 
    6.30537925211171, 6.56037541472346, 6.92962147972619, 7.33861622002132, 
    7.74016820390764, 8.00670798696016, 8.17043296298128, 8.16579113624364, 
    7.90400036604982, 7.57817182932429, 7.30559462992765, 7.09241328707552, 
    6.9283162237615, 6.77941805324977, 6.64082222429357, 6.68638739908077, 
    6.78289103694883, 6.85285794914596, 6.81013544690014, 6.63632776725734, 
    6.47595864898771, 6.39095933633339, 6.44511757908214, 6.57348502580371,
  7.509557889572, 7.60759308715627, 7.70343071772099, 7.77103341097608, 
    7.79351562876318, 7.78026829706714, 7.73612087956802, 7.67124253301731, 
    7.63472584018928, 7.62498796413439, 7.58648430617484, 7.49970262055789, 
    7.40422571820837, 7.37525736250822, 7.47993960085935, 7.68468190144245, 
    7.94283014244338, 8.197077159737, 8.46766983060778, 8.72948567222205, 
    8.953935880736, 9.13736773266626, 9.25756987731397, 9.24873197098894, 
    9.0883488514067, 8.8117594268852, 8.47933187387114, 8.13706178309774, 
    7.79345060530657, 7.4829539671479, 7.28820923964898, 7.23414932089519, 
    7.28368036043642, 7.38319881913399, 7.52834747118711, 7.77882021715849, 
    8.13018840766185, 8.49070670517961, 8.85517576025532, 9.19604173322008, 
    9.50313319014295, 9.68170308703106, 9.71028816845661, 9.59683804684811, 
    9.43839126828775, 9.31896045514755, 9.17410472878807, 8.96485843195867, 
    8.72664848524719, 8.4705121017175, 8.30092458128881, 8.21803000280567, 
    8.14714525585436, 8.03292744638349, 7.88026968731509, 7.76832308018413, 
    7.68129740309841, 7.57224839887039, 7.47512524756808, 7.45637223893865,
  8.6706529934956, 8.74896880864554, 8.80051272599741, 8.80942399261278, 
    8.79469875934741, 8.77926789655008, 8.78257071705114, 8.81633693471404, 
    8.86505495980976, 8.92190852489898, 8.99386465271147, 9.09575869254313, 
    9.24144925595653, 9.43513008022096, 9.68145300426693, 9.95601859142881, 
    10.2681728243827, 10.6043357318446, 10.9224212163659, 11.1866111811172, 
    11.3716688001508, 11.4356312881022, 11.3597486015129, 11.1498732875446, 
    10.830498920936, 10.4484514511215, 10.0422983037892, 9.64670457803505, 
    9.3137390835534, 9.11477579263893, 9.05521648198951, 9.07241213584753, 
    9.11947920471098, 9.19091338931741, 9.30122937989846, 9.46745581413675, 
    9.69612728610641, 9.97790779560253, 10.2920944624548, 10.6312948379973, 
    10.9453789387872, 11.1890085485949, 11.3519525018524, 11.4493068403774, 
    11.4896034634971, 11.4440888093533, 11.3056336318375, 11.1028878635373, 
    10.874350523678, 10.6504755090696, 10.4133732360225, 10.1267288911971, 
    9.80657581530086, 9.47354594766286, 9.16830239373206, 8.93356310257577, 
    8.75352871483313, 8.62669679379416, 8.57848419075832, 8.60152838534088,
  7.46032006482548, 7.7811957475718, 8.01453362201818, 8.10521813079334, 
    8.03256248667238, 7.79416990788803, 7.44751655223958, 7.13612448934124, 
    6.92624628624435, 6.84077529985551, 6.86015187799218, 6.96974081129566, 
    7.13559006001984, 7.32321684910993, 7.47451613944752, 7.5679427566472, 
    7.55149144457555, 7.45111707485437, 7.27567475323952, 6.99931322781209, 
    6.61369172783142, 6.15034653949557, 5.63710210386886, 5.07349481238706, 
    4.41544173776117, 3.67130358666982, 2.91542505642862, 2.17281972651171, 
    1.56029218554505, 1.10315367341363, 0.811898352773331, 0.73544418078278, 
    0.903414486707507, 1.29320589504599, 1.91144658591528, 2.75148076439673, 
    3.78145665458749, 4.92502186248109, 6.08189940075896, 7.1409199262677, 
    7.98125647973869, 8.52900418007565, 8.80233857173397, 8.8356416710589, 
    8.55505091345721, 7.9623722077806, 7.21807828540769, 6.49059089754846, 
    5.84885608119982, 5.33530021726567, 4.98276623441474, 4.80741097840022, 
    4.79691063433811, 4.9348176894668, 5.18273207003425, 5.51490396909663, 
    5.8870526946728, 6.27037554317184, 6.67531780002347, 7.08390782718818,
  9.94395920407263, 10.3762420288265, 10.1323838528778, 9.27234635259806, 
    8.1062515640512, 7.08741924354596, 6.51867207045124, 6.52549500013794, 
    7.20921342517116, 8.46832174521446, 10.0222696018612, 11.3960409146367, 
    12.2185301110899, 12.2704770727583, 11.7085469433899, 10.7286568256816, 
    9.78044839280477, 9.05206118984401, 8.86075853927829, 9.45365245677564, 
    10.4667017838707, 11.2471163639693, 11.3582317575107, 10.6502583819933, 
    9.19122996420024, 7.3479269528698, 5.54731485005255, 4.28195885510329, 
    3.61427200186311, 3.45531556024155, 3.66120434246694, 4.03746004983538, 
    4.26757143646489, 4.21030122286761, 3.95868678613485, 3.79836512890206, 
    3.97759358675691, 4.67572881168685, 5.92284282941042, 7.6088955238964, 
    9.46347344141615, 11.0617826648191, 11.9660562477514, 11.9623472018202, 
    11.0389410699922, 9.22640854609941, 6.9894157233909, 5.11562334393379, 
    4.16552210522432, 4.22973975861264, 5.02133499114069, 6.12686333791106, 
    7.1136769333944, 7.62064049798847, 7.54835118964919, 7.18853984093574, 
    7.02710879299095, 7.36822608160918, 8.12786690048994, 9.08739622454573,
  9.41766979402565, 6.95436141955774, 4.16636667524446, 1.86729061610868, 
    0.813428098628892, 1.32703799784976, 3.24786779394656, 6.00752671194281, 
    9.17632426560568, 12.435303485822, 15.4752696151095, 17.8552467544533, 
    19.0447574746822, 18.6487483607814, 16.2310998996, 12.7559415047662, 
    10.0350727932104, 9.76534292236367, 11.5194620789563, 13.6733189523158, 
    14.7498652008827, 14.854600047411, 14.7146236387184, 14.3097286045523, 
    13.4774506596144, 12.1025899649662, 10.3043832601334, 8.6767139258274, 
    8.39960792550468, 9.60662684187398, 10.6019956647629, 10.2554633910969, 
    9.08898830646603, 7.73047725801551, 6.70296773428196, 6.41387047132312, 
    6.99046412996743, 8.35468053679883, 10.1896540495006, 11.8346251063179, 
    12.6160602164181, 12.3600075103476, 10.984035675269, 8.69086995211214, 
    6.4030987658126, 4.97371519684567, 4.89132171466588, 6.37368215543997, 
    9.09818248160527, 12.5609591979278, 15.8748603308205, 17.7170770695771, 
    17.9477688500651, 16.9404092386133, 15.6380111642539, 14.1913523298935, 
    12.9283199600176, 11.9861777454388, 11.4937572578958, 10.9026737234729,
  10.8441928819411, 8.47512279457581, 7.48477809611061, 8.23696562875906, 
    7.32801177671892, 4.47055454253041, 3.08685628780025, 4.55611726457397, 
    7.34574612615691, 8.79677536302213, 8.30344557232877, 8.21543997531767, 
    10.4196647661834, 11.9774502010846, 8.70642810171028, 4.43181928977498, 
    4.0113672285054, 6.03720310643489, 8.74171944254234, 11.7640411423184, 
    13.8736937033471, 13.8402788731827, 13.2012746176514, 13.5169568413471, 
    13.3285920244648, 10.9876186926403, 9.08845658094866, 9.43307904798419, 
    9.52206977850343, 8.35828639935593, 7.79440676201288, 8.25614373595312, 
    9.18958986043388, 10.0587483598867, 10.1425803911141, 9.21385687621338, 
    8.75068375570834, 10.1288416863149, 11.7278305330214, 10.9728225313466, 
    8.50776878288477, 6.63783466278406, 5.50473708043411, 3.86597530228456, 
    2.84731573543261, 4.27475577671511, 7.38370888849393, 9.31973490531011, 
    8.57512085664771, 6.59321905877858, 6.82849831511474, 9.22005055599112, 
    11.7597468983503, 12.3698363555652, 11.3964813086043, 10.2012203572136, 
    8.24143537205073, 7.00949549925352, 8.58694947876991, 11.0784225520912,
  0.542658217385209, 0.989526842833734, 1.03897386620263, 1.22091370834626, 
    1.32510651744513, 1.85681001589877, 2.68811003108278, 1.2383974611535, 
    -1.49605328366172, -3.025452999123, -4.29678543950328, -3.38258617460962, 
    0.348425738722769, 0.951932644960811, -1.63560354057049, 
    -1.89548339899975, -1.61527607074574, 0.219101122003608, 2.8091568051021, 
    4.36795539506772, 2.94085303014843, 3.02449257430661, 3.54775210685792, 
    3.66494681066266, 4.61333239676956, 6.33228583506237, 5.81672496701169, 
    3.48955329545695, 1.04136910507165, 2.94356180618071, 11.2546287139008, 
    18.1453072806427, 19.3739041460368, 17.6290037793953, 14.9855948527951, 
    10.9670129624136, 6.99141339846696, 5.10458725760012, 4.58448469787329, 
    3.71959081436976, 2.17776171999278, 0.0692326054182461, 
    -1.53231039960639, -1.22996173051968, 0.979916759613324, 
    3.27789096595259, 4.20388812886025, 3.14955901087773, 1.11049505229917, 
    1.53994238429714, 4.28753447971491, 4.67046063912275, 3.79851832957498, 
    2.06648039429126, 0.479318632765679, 1.4857018896749, 4.37224409686571, 
    6.26057526942715, 4.26767074470666, 1.11328845591281,
  1.85197408073932, 2.91793650410486, 2.82980107033619, 2.78970330122301, 
    4.78835089618533, 5.70403792135108, 3.76584991831077, 2.3980482240022, 
    1.61423387598158, 0.475559746554913, -0.817796577126047, 
    -3.04271316299998, -3.89804907802125, 2.67518247164008, 4.29811873040698, 
    -0.336931892021859, -0.0503949615644375, 2.24180122618018, 
    3.78575450396266, 1.01890235927629, 0.49826421087458, 0.736830061016143, 
    -1.28759107166065, -1.65720829271206, -1.5372956266673, 
    -1.77489151195431, -1.86807703922437, -1.64891198915641, 
    0.93632538002145, 7.4028066831697, 11.2473517777313, 11.3360535889416, 
    8.29834080930684, 2.86489794342699, 0.675048643330465, 0.210545366610806, 
    0.0673439220605969, 0.321893506513124, 0.605227832453096, 
    1.75726037296024, 2.98625105286238, 3.06791237800101, 2.94495552704432, 
    3.54544861058771, 5.56292535783778, 8.28501987783606, 10.7569627953477, 
    13.2389806950377, 14.1951221969005, 9.48664488481779, 0.97685443154348, 
    -2.92359312713977, 0.306673293246132, 0.438681288179062, 
    -4.55126063353067, -7.88974997089849, -9.48348215312441, 
    -8.63995806070735, -5.01617205318284, -0.817878573980001,
  8.34141734549845, 12.1881589903371, 13.9576603893985, 13.1009995314401, 
    13.2733020283473, 15.1307853590139, 15.8881695107357, 13.9613802493611, 
    10.6207410549225, 9.12423140287186, 10.4652015952127, 12.1546970351928, 
    7.11668462199138, 0.420844367626715, 9.64076654782563, 16.9753884390765, 
    9.3499159302225, -0.135240333217082, -5.07441227144452, 
    -3.39417349119434, 0.337438668381067, 5.74380559906632, 8.55820863229203, 
    5.76921505329021, 3.16223083901697, 4.09037811897574, 8.1266780442301, 
    12.2384987403976, 13.401642604002, 7.71506192009308, -0.621106001222846, 
    -2.1619256619229, 2.19302238349403, 6.21091786508224, 9.92951186079073, 
    14.8656631829348, 16.5348954853957, 12.2420263038323, 6.02078448453753, 
    3.54041035963483, 6.17507820920264, 9.81683679318941, 11.798707193779, 
    12.6474044938995, 11.5245859723969, 8.66580664621712, 6.03003158514791, 
    5.74337449259637, 10.1442697724801, 15.4030111923235, 15.5762544568325, 
    10.5825254073196, 5.14270143732227, 10.2230072359957, 15.7285566476991, 
    12.7926309829551, 8.14316758750626, 4.82558143089615, 4.38604548153179, 
    5.57697707765429,
  18.4600928242134, 23.4358841939674, 22.899779726091, 18.6247455068742, 
    15.3881762576728, 15.2406250565628, 17.6124097545232, 20.9439854405787, 
    21.8267824738223, 19.77269537719, 17.2769136900664, 16.5327304030645, 
    18.7665271239201, 16.6062972039119, 7.85241118008373, 13.3613562691617, 
    21.6982155086453, 15.5459395613723, 9.09239981351325, 5.99501382461836, 
    3.59917514689229, 4.73142939134823, 11.1186833232041, 16.2749609699232, 
    15.5637131954385, 11.8282126981356, 12.0178320960137, 17.6172639207817, 
    22.3878331067405, 26.0645056502004, 24.1358382879913, 14.6258015451377, 
    5.68804186068436, 4.51381353791535, 9.13670897384936, 13.7364119202773, 
    18.9103892882513, 22.421853231993, 20.0252165106399, 14.7202871270088, 
    11.11236498953, 13.050643188365, 16.6019512277103, 15.2503762013566, 
    11.9918481806596, 9.18689374466345, 8.32686148652646, 8.84017618428388, 
    8.12712808808241, 12.1564546855153, 16.477598307648, 15.5106082916264, 
    14.462040194582, 12.4001749387512, 19.8698472851526, 28.8959455252911, 
    27.1288156689326, 21.531124333412, 15.1746141389809, 13.1626981464701,
  22.7418308238768, 26.2153593007549, 27.9286960387323, 21.9629870660217, 
    17.5788656641422, 22.1532596713646, 22.3032191062655, 22.4400964466774, 
    23.8956761708554, 20.3845783916939, 21.7672141294678, 22.8880637367611, 
    20.6166551680027, 20.5666567059177, 21.7668530496128, 19.389844957053, 
    20.5181696447479, 23.092017056169, 21.0479764071045, 18.7988085883783, 
    22.545753492626, 26.0894078244413, 24.6102096218755, 20.7548881502578, 
    14.9512405559088, 10.3325821192315, 10.4387621695149, 19.7444601773694, 
    30.6139681772627, 32.328375557332, 28.287114708936, 22.4604797183981, 
    17.6076860611692, 18.1613372800638, 20.4102050829978, 21.9778029492437, 
    21.8944311364135, 21.1663037587209, 20.0959384780836, 17.3538727471908, 
    15.6532375103141, 17.275794086601, 22.5058686184013, 26.4908407820866, 
    22.8441121144372, 17.3744549801143, 17.9019958924257, 21.7596979227153, 
    23.0590363769884, 20.4040953488322, 19.7472036075113, 17.0527886111249, 
    12.9166949915288, 16.8835199450054, 21.793034027236, 27.8870410719039, 
    30.9748890034252, 23.1664582424289, 18.6298297316687, 20.5444473550245,
  29.7403280500383, 30.2678581345995, 30.3488417153743, 25.1374546712608, 
    23.7123762950174, 25.3921721856588, 29.5218777790277, 31.1769982790512, 
    27.1457422028559, 26.6357706037197, 25.4847825208904, 26.2799362301494, 
    27.6110711844032, 29.5289650570914, 30.2947297688544, 28.0115322996739, 
    25.7477358645225, 26.3687254693802, 27.2384186684187, 30.6502375552847, 
    33.810885160901, 38.0339634737107, 39.7092584287227, 31.8048741531118, 
    24.9512354654336, 22.4680340782109, 25.7179912456049, 32.3455145717248, 
    36.1474318738597, 37.8437877939044, 34.552105012529, 29.3898934375144, 
    27.7458070760414, 25.4671911495896, 25.5923833954154, 28.5945523841606, 
    29.3375377382681, 27.6825946558018, 22.3803188044658, 19.861682712291, 
    24.9158959217702, 29.9348858898786, 33.2734216004392, 32.9609156404378, 
    27.7679953161546, 25.6525018523958, 25.6061108752561, 26.0094338152101, 
    24.5945078759439, 24.6843799035666, 24.1437679386865, 20.3533873418789, 
    19.0194085898456, 22.7122766408721, 28.9438519223759, 32.3056994576162, 
    29.7734332719046, 23.440602917102, 20.8061762322966, 24.423703360338,
  26.3584611390548, 26.0303269071236, 19.0571906108014, 19.8633068266407, 
    21.4961239564224, 23.3279129357552, 24.9839928309271, 22.8221699144133, 
    22.7884046514082, 20.8308855525027, 21.9307818006372, 25.5393343393734, 
    29.4630952925935, 33.0371723503176, 25.3906720015684, 18.071379468368, 
    18.5050618936507, 18.5413134501992, 22.6718669125271, 36.3021296208624, 
    39.7307222899785, 32.3793292643008, 23.3519489340416, 19.8685505057445, 
    22.5274793731617, 24.0041941389947, 30.8203033523165, 32.0171475050105, 
    27.7367363501524, 20.4505013542446, 19.852238678324, 20.6353344992374, 
    19.8222932469811, 25.6207693589213, 26.8849741152769, 26.4908511072091, 
    29.8787564954082, 25.2909342242536, 19.2430921185201, 21.0451493675641, 
    22.0941507459799, 27.1663432878063, 27.7615174466947, 22.7101308161565, 
    22.6568350955654, 26.0283769015712, 32.3799107509385, 29.7014164204491, 
    28.9248343478381, 28.9699736066052, 24.364917657043, 24.3413268444983, 
    23.8914454386404, 26.3690708299056, 29.475959567723, 24.6863849827808, 
    16.9921369014645, 14.7232922795675, 20.3661173180102, 26.0839165026817,
  24.3047336883557, 17.2614972660982, 15.5982244516428, 17.1974360940862, 
    21.6163183056674, 19.9756068376027, 19.1890422127551, 21.00964810371, 
    13.5091202387714, 14.9072357416569, 24.4364731929668, 24.4135679735262, 
    12.8345478201372, 15.2472014008234, 17.2172558577606, 14.7551486500804, 
    8.63303168719467, 16.295855146586, 33.0793767764932, 29.4355541509751, 
    18.143587816586, 12.2979842538694, 14.7630600078577, 18.6196141201267, 
    19.3047680433028, 25.7594545896149, 31.679124518081, 22.7650775106362, 
    10.5342229076775, 5.29743098907665, 6.44183047825466, 13.4248018886983, 
    26.1827105330001, 30.1166219772615, 19.0792057528724, 12.966794188914, 
    11.8914803045939, 17.5893353294691, 19.1762161725333, 17.81652743338, 
    23.6685765696591, 21.1481688244721, 13.6616759884436, 9.51435211196435, 
    15.6837180761705, 25.9743919936465, 28.7090935623505, 23.1913076572921, 
    16.4896338904192, 16.4579983874339, 13.9649141051647, 14.7857602902669, 
    20.6807196179309, 21.7771945536631, 13.1096554784998, 11.8926243349359, 
    11.6284191233762, 20.2184027190172, 26.4106721641916, 29.4719339448091,
  15.9406034958849, 15.0553378079401, 10.5832811236704, 13.9513820493438, 
    13.5656091487538, 17.6835731707763, 18.4373148162397, 19.0833882358082, 
    19.8746019592816, 15.8877709965571, 15.5412764175355, 12.437549172559, 
    9.47032044738181, 7.82461141934991, 8.57017888070003, 7.26591446470335, 
    22.5680634961474, 28.813357467339, 24.099824712708, 18.4742943896322, 
    8.3245081141685, 3.34485748939542, 11.3280461148817, 14.6143243964292, 
    21.0889025429132, 17.9264762431872, 17.8721543402181, 15.0471954623654, 
    9.64455723355143, 7.39417767896031, 10.8799677310777, 12.9102720957569, 
    9.56028644950971, 11.4382129300924, 12.1419679311981, 10.883759391602, 
    11.2120776475474, 15.3498599114823, 22.8225222155165, 30.2697731751458, 
    21.7441304371135, 16.9063349674227, 15.8308972294128, 18.2376118921988, 
    17.469897031911, 11.0518973323546, 9.84421548284088, 12.2804880686608, 
    14.0001728295987, 15.819300294303, 18.1479221676344, 19.4087337305839, 
    13.3103491480115, 13.5682789392323, 14.3589638392017, 12.1311060851554, 
    17.9018628508359, 22.0648754934038, 19.5927158023723, 16.3587401910094,
  7.74899923151378, 8.95553198091222, 13.0379255038855, 10.6498840205712, 
    7.46985213315467, -1.8707582444566, 7.17757693694491, 8.267761618607, 
    11.8231692806787, 12.0406839296746, 7.13140658279225, 4.68429865917532, 
    5.00011540696198, 6.81299387232489, 11.8103549806982, 18.7053136528061, 
    13.0832819540286, 9.86343968246365, 7.03583189084068, 2.86836451353293, 
    5.02752313708704, 2.6455226071757, 8.19897092838733, 10.686842019527, 
    11.5880458284383, 9.99087137080039, 4.44443224132288, 3.61792279336627, 
    5.6725178219685, 8.75538229883219, 9.41358071819204, 8.60861631410006, 
    7.80268453718326, 7.48135847027291, 9.64491808633469, 10.7622462158429, 
    10.7132926771086, 9.08125114724586, 5.57752730840391, 3.53082013551667, 
    7.08227849387377, 8.86393410158876, 8.80393543709758, 9.97442543572839, 
    10.6895446587103, 9.36877410617187, 8.03249031354213, 6.09776991460339, 
    7.244481739807, 9.84965747955635, 8.97514066995189, 5.86880328494157, 
    6.81299342981445, 5.49865675541359, 7.24825664197541, 9.96662047645944, 
    7.50262493596714, 9.26410369825448, 4.62078240078134, 4.66465521150385,
  4.6443473477012, 5.76216566577162, 8.13944969683475, 9.90018585645157, 
    3.45296067533812, 5.27591648816218, -5.20594056171316, 0.677602890702147, 
    5.37983263445271, 2.93590186381158, 2.8018153273417, 6.11307756946892, 
    9.29030180778665, 12.1159021329078, 12.5664917918168, 8.99976835376141, 
    5.00979809314441, 7.78164762698346, 6.88981989814563, 0.443855101638615, 
    0.840045400809784, 7.59175254803446, 7.63349054286074, 7.84026384629833, 
    2.9416709779599, 1.72494590681503, 2.81999162734167, -0.537007617522777, 
    1.39981580255997, 2.19078074989504, 5.28092722959861, 9.32616286798764, 
    8.74670760627239, 5.11879932075951, 3.53427628500029, 4.22714333740927, 
    3.70251969518646, 1.65312834914508, 1.25502615857227, 0.0476125276479502, 
    1.68853599288525, 1.18038232707092, 0.930961300686657, 2.2676018737881, 
    1.4804799403949, 0.645688377468891, 1.33386645820049, 3.10260771234706, 
    2.02035299601399, -1.29374601439398, 1.51434470020111, 1.49257110470745, 
    -1.5733058573459, -0.285093969003451, -0.436809115258874, 
    3.18009508519678, 2.00630073397907, 1.46812255812353, 8.91015534792611, 
    4.06409017571534,
  15.5636244321971, 12.0975660231522, 12.3646812608663, 9.49672636391409, 
    8.16070451635095, 9.56493775818846, 3.38176368150906, 2.20686494673111, 
    11.1222362067603, 16.6926216091347, 10.8229847396463, 11.2511539608766, 
    13.3779801563622, 11.3602143341857, 10.0187159104193, 9.8378270305015, 
    8.55243898183857, 8.8577747661515, 7.26890415110069, 8.74532884528631, 
    10.1372166022478, 12.5545880586371, 13.1444664965924, 9.47780573495634, 
    2.72810061876104, 2.33702194577593, 1.66290838820877, 2.16216709355974, 
    7.90471437077203, 11.9796547977044, 10.3489146019316, 6.30113015056514, 
    4.61694455897083, 4.35366259402109, 5.67816601932716, 8.022236807395, 
    9.40733582098802, 10.3354885463354, 8.89968094130329, 8.61252155377654, 
    4.75057222267305, 1.85626093746542, 1.5739667694887, 2.86529289012529, 
    5.91446100682335, 9.2165239581165, 10.8446873711122, 8.71914017601901, 
    5.2253827376838, 1.3817693271465, 4.40880850629966, 4.77680077191135, 
    5.69383187525193, 3.16265903525555, 4.06191466530535, 2.89459652076495, 
    7.42411440704114, 7.37653725272247, 17.0665371519742, 16.0666028124525,
  5.31690760045402, 13.5922239647196, 17.1957448934295, 16.561621551121, 
    16.877777300136, 16.4546047144764, 17.5161267265634, 18.5944792852159, 
    21.2917376093599, 28.6271346488243, 26.0441824241927, 18.3174073163656, 
    15.9860547428513, 18.6316271122305, 18.1297841495724, 16.1268173357856, 
    15.6200134491727, 15.1038021467631, 16.3265357612338, 14.9499763057148, 
    13.7911774606811, 12.3722058131143, 15.2502449253958, 19.3674137627351, 
    13.3526188292514, 6.5547035365793, 7.99764331802183, 14.5889163062132, 
    18.9027048650225, 15.967753193527, 21.6548008417196, 25.7116032114339, 
    21.618258358371, 15.59426098067, 10.8168622279959, 8.9380403465535, 
    11.0520843511081, 16.1619819817897, 23.0791830870985, 22.6309098188981, 
    18.7759249905414, 15.3971511264612, 12.6289007552886, 10.507614614476, 
    11.1653892869861, 14.3875239945428, 15.8082679054358, 15.3332863434134, 
    16.1062054191065, 16.8268491695236, 17.3988762086824, 16.4793761837277, 
    15.6689304083597, 17.6662779049288, 18.3418890356907, 16.3688980238175, 
    13.3196183834768, 13.4995159226405, 17.2603192394622, 16.3653579473353,
  8.18925292727205, 9.41977311292309, 15.1536165736821, 15.6783599294132, 
    12.0442773445061, 14.2775451711036, 18.3026735160392, 19.7458011282885, 
    23.5036242579341, 25.1248955094894, 24.1138172019408, 19.0015787464136, 
    9.47853987531153, 11.3388974467067, 20.1539129900504, 20.5804130428667, 
    16.4173453034317, 15.7017792411464, 16.4480754611525, 21.8218409634742, 
    19.1558570981007, 15.2503273938255, 12.6221969811686, 14.0584941343942, 
    20.3987452189042, 23.2509567884541, 21.9028655870296, 20.4144239565755, 
    23.7907486146075, 27.8499090142454, 20.7399145804984, 18.6525285097113, 
    22.8541830312545, 17.3581739263962, 11.1929643500001, 7.33980207646699, 
    7.8419179584021, 12.8261246478649, 18.819880817364, 25.654255788601, 
    26.1335827865438, 17.4734453074468, 14.3854784993956, 16.8221593332414, 
    19.2239970674161, 17.1592073280283, 19.111757825037, 20.5256800207297, 
    21.0587153532882, 24.7643809265335, 18.6351310357213, 11.6582408516633, 
    9.93585557524244, 9.05284488551389, 10.1507927398551, 19.2145621287034, 
    29.3160638739725, 29.3485981096466, 29.599726295236, 25.2904781034927,
  24.8717254381435, 24.2186843564604, 21.1860059409163, 20.8684507971413, 
    18.2293185181806, 15.132500684795, 12.0216089100174, 9.1698392834831, 
    10.3320599873302, 15.3251620653561, 22.6501637984077, 24.1853932794976, 
    15.1080118385417, 8.34099365739866, 9.72143691193152, 20.8098797074174, 
    31.0341916791533, 27.5258362902166, 18.2806884613966, 12.6882454527943, 
    17.0213218363807, 23.8889101728919, 22.5562397871989, 18.6125858953644, 
    15.4757576039179, 17.6497118965516, 22.8896483346676, 23.7326933827499, 
    24.4699551235068, 21.6318038575681, 23.0302429350116, 21.234657521592, 
    23.4008396992747, 27.3813997128027, 17.6365147359534, 6.83506890944063, 
    6.1067663116052, 9.09024718050372, 13.621548368274, 16.0672997011662, 
    19.8426616733353, 24.8237578286919, 22.7313821302079, 16.4212823717787, 
    13.5202837809149, 12.5640165323467, 9.98775642511833, 16.8830499662226, 
    28.4859899739146, 25.5827781082546, 25.1876794125987, 26.7748985538104, 
    17.5109063778644, 13.8062679419115, 14.6099878535424, 19.581608034006, 
    17.5729099858332, 20.1590925764114, 29.3060511933769, 30.1089215384785,
  32.1982708780704, 32.5724831112834, 27.992658522801, 23.0312658320671, 
    23.573715800529, 21.1347689887344, 20.0007312994937, 22.6589545074099, 
    23.8711669757748, 22.9068130864795, 23.1448892924946, 24.8389980603744, 
    23.8719846107334, 17.9125438015671, 16.0142007889951, 19.7828174203748, 
    25.1094569196492, 28.7270840023405, 24.6037638421932, 22.914061530747, 
    25.1537326388519, 21.6683737166375, 19.7854792292849, 25.28127131794, 
    31.0626011296703, 27.8705236768931, 22.7423620583038, 22.1124962320469, 
    23.0538300821425, 23.1889688164139, 21.6279847519849, 22.2355300591916, 
    24.8764039943679, 28.2625476485922, 30.1146183091947, 30.4669332926245, 
    28.2213248985397, 23.9445386479895, 21.2422549279085, 20.6876295536747, 
    21.9909619232876, 25.9142143421402, 29.0961649725145, 27.5098761500145, 
    23.3714884479648, 23.3266755765774, 25.9985494307982, 22.3934841317987, 
    23.5155954441747, 30.5283235139179, 28.9504594793016, 28.6159474691586, 
    32.0855386047297, 32.2230978981931, 31.7338825839326, 29.0555744799275, 
    28.3977782978207, 25.3982901779352, 24.4232769187384, 30.2209728696588,
  28.0284287742178, 28.7102857740519, 26.9672447774424, 26.4162302126503, 
    28.60788950328, 34.2411028064441, 37.2112643270967, 31.9265898231963, 
    23.0011116931109, 16.6789426188434, 15.4380692207213, 18.3144346513694, 
    23.3840410140622, 27.2140806299241, 27.0170688791059, 22.6419772046755, 
    20.2449590703474, 21.6117367485471, 24.9475169406308, 28.0033759383417, 
    28.2015104967153, 27.4230519994404, 23.4148053147156, 20.7047145865056, 
    25.7992927401378, 27.4567129029888, 22.5110327887734, 20.5261723886462, 
    19.2783053777486, 21.2000020826711, 24.7632383430974, 23.9513179048171, 
    22.1009908911784, 24.9309148496354, 30.8734322493857, 32.8456698242824, 
    32.2325238264325, 28.9840688762973, 22.4221733537134, 17.1661018166185, 
    17.7293639998994, 20.7542373867981, 22.7358244853491, 25.0321851936556, 
    26.4685736789794, 25.5561917752943, 23.600491894983, 22.4725441514071, 
    23.2682942646832, 26.8514390931492, 29.6986924227764, 30.3736426257757, 
    30.4193474624174, 29.1904021938928, 27.4393642499497, 25.2257403273876, 
    15.9580513174772, 10.996190399416, 12.8512629958394, 20.122388885898,
  24.7841053212643, 21.8607060376705, 16.2331591583445, 14.2569645456331, 
    16.4980361495933, 17.893794776452, 18.8684825713536, 22.0734827384192, 
    20.2876254291301, 12.9582495190727, 8.21491915102379, 12.5491323425873, 
    19.9303564333177, 24.7913466859061, 25.9201422815639, 18.821828741837, 
    11.9235785107485, 11.540979555719, 15.7207561211807, 19.0875847755504, 
    20.6773590738264, 21.206429320712, 18.1829850095861, 17.5218717218706, 
    14.3045692215167, 11.3494746175523, 13.5315436178034, 12.347783090415, 
    13.3313194780109, 15.9541154643477, 14.3643079573928, 12.2214551824275, 
    10.408665970838, 10.1301804766895, 12.2229014495284, 19.1976232683572, 
    27.7837910030374, 27.0395132295794, 18.5675955296606, 11.680017009726, 
    8.53437136217699, 10.5381490458389, 15.4536917396135, 16.8006877226923, 
    17.7894384465048, 19.1591280403857, 17.2998942215629, 16.6808528918959, 
    18.4597372652996, 19.6558128592282, 19.6828104569477, 20.0604080895894, 
    22.7377961244682, 26.0417097698029, 20.4007369546388, 11.732903711672, 
    11.5621111287082, 13.5147248352347, 16.9147478028307, 22.4390315440702,
  -1.77370688047216, -2.13121831883207, 3.3531753359068, 3.95149478211949, 
    3.91297040489927, 11.6443708677447, 22.714872207744, 22.5230333270132, 
    12.7677447717385, 6.13959658091099, 5.5745917483993, 9.72701689624653, 
    16.3066429719613, 19.3790225796369, 18.3798128568879, 17.1027843722366, 
    15.3122145120289, 14.2041089573759, 13.3900498779809, 16.2847889577543, 
    22.0448792459239, 18.8663020100703, 7.42522308763775, -0.580574225908062, 
    1.07744552799621, 10.477864778835, 14.8513618828764, 14.8448739254591, 
    14.1054552230484, 10.4700666871331, 6.46941037856519, 4.71311779747177, 
    4.38762998768798, 6.25544668118914, 13.4781245808345, 22.5541681192905, 
    25.3787773004247, 20.2693814558112, 13.845607243234, 9.4686995267715, 
    8.51852507203835, 7.5390422648749, 5.13945135102116, 9.5581559151021, 
    16.5724401620134, 17.2343452728693, 14.2034593826687, 8.52166354755022, 
    1.82607020053699, -0.259577840244494, 1.03807087985145, 1.7700922764764, 
    1.04206662613249, 0.598722643000237, 5.55706670454382, 11.8433077509343, 
    13.1446323647135, 10.5759374990506, 7.68859051589409, 4.6360259717621,
  5.28456851851909, 6.44263083052269, 5.23808072869502, 6.49899526365623, 
    10.1086242426842, 11.5093480372581, 7.11565986393291, 2.57264033873026, 
    2.69743320634159, 3.99222340059229, 5.40449025814326, 8.30778062891035, 
    10.1495831726125, 10.8985031049174, 11.3062106574208, 10.4174093893527, 
    9.61470576714367, 9.41123294330475, 8.82909400552671, 6.1301916521626, 
    -0.755359305108151, -4.83203218213094, 0.0548644915289781, 
    5.43663073583854, 7.55863715812078, 8.42038029437956, 9.28902243158512, 
    10.8661256896999, 9.64468360465908, 7.78785497873513, 7.17389027312391, 
    4.29354792097133, 2.3913689406397, 5.82280656387315, 10.0704475754538, 
    10.6862246114089, 10.0350998969006, 10.0554947399623, 10.205321567285, 
    9.70073068096051, 6.62558679818544, 4.62013125311152, 8.21669519032363, 
    11.890308185506, 10.7343680185243, 5.78629845948228, -2.46732330513093, 
    -8.45517272647207, -3.77073611123083, 1.02230561257412, 2.4732156984479, 
    3.58245061478666, 4.2657265421078, 8.95450722521373, 13.7251131373098, 
    15.1999612408263, 12.7173009824988, 7.38079184742467, 4.62095124643486, 
    3.99945212793176,
  3.80845976218267, 6.91937030799558, 5.59909240916989, 3.52262173043492, 
    3.61462704714915, 4.33267376479288, 5.17488615801741, 5.62442961110805, 
    5.79063187257492, 5.63798691791854, 4.81094100422938, 5.0563911442345, 
    5.35702540512, 4.1983590708827, 2.36527086865126, 1.0649646542462, 
    -0.0560698802267546, -0.540042328865169, 0.199606965983521, 
    0.231278395530141, -0.56652603469788, 1.14806440290455, 2.9685202468504, 
    2.66132227699168, 2.55500859141355, 3.24774114114924, 4.05849023463341, 
    4.34397974208024, 4.55596003389037, 5.34192113441735, 6.62725298764744, 
    9.82162139268141, 13.1051383343262, 11.6012606730114, 7.59780527645852, 
    5.44570018512858, 3.2920648176157, -1.26367657655637, -4.66657886841729, 
    -6.31486323200169, -4.96645114572039, -2.38453961217459, 
    -2.32044706696845, -4.43900704380973, -6.03792450733794, 
    -3.68042182334517, 2.7023906031096, 9.72391719847607, 9.7983845288427, 
    1.75668314821155, -0.952951525899087, 3.80823258280608, 8.437256620217, 
    9.06416751253974, 7.90564284901847, 7.97556673708921, 9.05352793104886, 
    9.16346938834724, 5.84512565994504, 2.71088314256765,
  9.49146170599055, 10.0873214310928, 9.30708248634251, 7.89028335633684, 
    7.50672667648866, 7.49200543890802, 6.42620203867221, 5.99813224017419, 
    8.00350749418223, 11.2539008220994, 12.3253477611316, 10.1938575008796, 
    7.04718467633103, 4.81107166758108, 3.09245602075081, 0.429670820874296, 
    -2.34180662488088, -3.56549757331872, -3.0241888586881, 
    -0.781975651711003, 1.82557234156972, 3.32890198186232, 3.03632428500545, 
    1.51113881613532, -0.0289425312232899, -0.709157711844655, 
    -0.46824529620541, 0.345266093861246, 1.42519158790638, 2.93232521978322, 
    5.02719346468191, 6.84866885504155, 7.51981676429961, 7.23106705755664, 
    6.64643237869411, 5.41253014562193, 3.7472458926404, 3.10691200856596, 
    3.97713335358449, 5.06462092332465, 5.48772062973683, 5.60458316117661, 
    3.54349744750447, 1.5581521020817, 1.18054789109296, 0.141924378093491, 
    -0.665209436592056, 0.976776550224065, 5.08846346953842, 
    8.35873540099231, 7.13826514866183, 3.38409255224008, 1.6136485285521, 
    2.12154607052361, 3.83456254593734, 5.76809983213974, 6.9073822245221, 
    7.27677622721947, 7.41156700166545, 8.30260900364248,
  8.09579110868516, 10.8715414186509, 12.5464045371733, 12.7597376157071, 
    11.7398384673092, 10.0723784005292, 8.34950082551, 6.98818077502934, 
    6.52116897901786, 7.33666856693285, 9.28605577747615, 11.4840603257584, 
    12.7232876416234, 12.2600372687192, 10.4966979656047, 8.77008536470827, 
    8.06514424723465, 8.17875853558597, 8.02200940721717, 7.44033469795326, 
    6.44470086992806, 5.52970627573591, 5.11785011599992, 5.4762357005629, 
    6.33667372660451, 6.87861645985787, 6.39317568337907, 5.15626242525821, 
    4.30791942406985, 4.3265887509267, 4.69267464015534, 4.9575955862517, 
    5.16797812686289, 5.44475469234386, 5.35573743033676, 4.40306205703329, 
    3.13044110827267, 2.87116527275979, 4.78386468497969, 9.09877410325183, 
    14.0284545283203, 18.1793732082354, 20.5777696907835, 20.8498966050404, 
    19.2822888841352, 16.823548082971, 14.445723244241, 12.3403848653081, 
    10.6830892934981, 9.52453043666803, 8.20756744595032, 6.37594339652559, 
    4.47373839128816, 3.13269657944033, 2.55918324881671, 2.46653752377491, 
    2.410245806554, 2.5220134784602, 3.29276625814784, 5.23209858130399,
  4.88386630607035, 5.69777741332706, 7.04821357288923, 8.4583016759482, 
    9.37592189989038, 9.45603897078762, 8.65520171534667, 7.32978040094754, 
    6.04892402168341, 5.2933179786687, 5.1935298794413, 5.50736346992968, 
    5.84316472484015, 5.99882581372876, 5.97334624242615, 6.11793538250476, 
    6.65861792722298, 7.89178511353348, 9.77309005513579, 11.8452164941844, 
    13.7271019930637, 15.1378496601991, 15.9722507759552, 16.2734093330125, 
    16.062217371961, 15.3868464758152, 14.2970078487433, 12.6952528121698, 
    10.6220751162282, 8.31529818959301, 6.30696815999639, 5.18148553917582, 
    5.24439083137204, 6.37231072907056, 8.08644328647188, 9.72295599465018, 
    10.8655866200071, 11.5852268403473, 11.9195712190159, 12.1062342387432, 
    12.6876265331173, 13.5766831786845, 14.2777771216156, 14.3968817342524, 
    13.7894929320324, 12.6365781559117, 11.2229706307624, 9.8388600214179, 
    8.72122922576649, 8.08668003701963, 8.04328071107294, 8.5246930833398, 
    9.24713499255837, 9.76972013992273, 9.73361195370164, 9.03494477696022, 
    7.93014280202802, 6.70449154501063, 5.56584007325851, 4.85138581216761,
  4.14002315170251, 3.67200544837813, 3.35693969569962, 3.18073560915184, 
    3.10464953519041, 3.07992036031573, 3.10504628828086, 3.19514012924289, 
    3.33908406205257, 3.51365379542359, 3.71834688011904, 3.97378838975479, 
    4.3026630723953, 4.70183408333204, 5.17954973399003, 5.74937579257756, 
    6.38500846712922, 7.09030614474046, 7.87026928243053, 8.75057280148524, 
    9.68592382772715, 10.6043789971071, 11.3840364777882, 11.9395809280575, 
    12.160755604566, 11.9641454321368, 11.3660289465913, 10.4079889548755, 
    9.1193506962305, 7.68758923246338, 6.31746587143658, 5.15920025762625, 
    4.27543570360979, 3.68732181830314, 3.37600644709533, 3.29975655666797, 
    3.41090000318412, 3.65826429422876, 4.00485621178216, 4.436438960569, 
    4.8910648761201, 5.34195521995465, 5.80825821046543, 6.28285329915873, 
    6.73893438898442, 7.14149225594289, 7.48266119989458, 7.75156707000631, 
    7.95229971189747, 8.11102443085896, 8.24069260748904, 8.31990674049873, 
    8.29765891754506, 8.15174716283569, 7.85140888418772, 7.36519830336645, 
    6.7777693687357, 6.13393012617851, 5.42043501411828, 4.73225835261593,
  0.420392587166876, 0.927116837020153, 1.50287095630537, 2.09519138608497, 
    2.63031131386266, 3.06781563444745, 3.38336521981497, 3.61926838395001, 
    3.79908370327612, 3.93026927759214, 4.00708618309716, 4.07042708248612, 
    4.13987240187512, 4.21923868647483, 4.31701500931243, 4.41660555948528, 
    4.4596058601611, 4.43422861371976, 4.28477698098604, 4.0008913949285, 
    3.56879476753621, 2.9766921872527, 2.31148436406648, 1.63059158349914, 
    0.938328032433093, 0.190031861463878, -0.535277485188578, 
    -1.10384651739857, -1.49213683679162, -1.69568336886059, 
    -1.68779912783382, -1.5285484907333, -1.26374107087879, 
    -0.917045270787188, -0.514260792350932, -0.0864253051558309, 
    0.371839634302359, 0.877746503204203, 1.4241677828484, 2.01043409514731, 
    2.60567175543004, 3.14499580876977, 3.58243858934845, 3.96928785164779, 
    4.26231690887292, 4.31175196778536, 4.12978639076369, 3.82879539502771, 
    3.43083481860292, 2.9279406738143, 2.34193650262641, 1.7316516768074, 
    1.1558551466378, 0.638643495369485, 0.216445844736023, 
    -0.0941705632709402, -0.286112031430207, -0.330081878226132, 
    -0.220740876625558, 0.0345041047896912,
  10.7491698276962, 11.6933481410354, 11.9748866817596, 11.3944138176626, 
    10.0982746930453, 8.45109919680755, 6.90961470456984, 5.70223884570904, 
    5.05145964346004, 5.15034747528692, 5.98220044656112, 7.11916349681004, 
    8.01904072671239, 8.31938088838656, 8.02460141490422, 7.37657004149148, 
    6.72520046883037, 6.32158983540668, 6.07304767603834, 6.44685314762508, 
    7.28652956573018, 8.00031961664602, 8.20394038832838, 7.68710469826738, 
    6.34567181235378, 4.52260228284723, 2.75060662071319, 1.54861895212523, 
    1.16887611920035, 1.38112638067093, 1.68619370230737, 1.78310304665542, 
    1.52287493489284, 0.869329856866318, -0.0234423013967634, 
    -0.765007705905197, -0.997258923089128, -0.452387247058729, 
    0.988536029723602, 3.23517296154228, 5.85786503485689, 8.25330935795549, 
    9.8653156304773, 10.4270991807886, 10.0397956125707, 8.71278504521783, 
    6.52799350856468, 4.04952432899257, 2.01585578566608, 0.877675182197924, 
    0.714719637247772, 1.27660885102488, 2.20061287752523, 3.13532131812032, 
    3.86374062912797, 4.49597541624304, 5.31397727052311, 6.45990272975331, 
    7.86263235539974, 9.37620580503356,
  7.03377079680545, 3.96941941659418, 0.622797033020705, -1.6094191250967, 
    -2.41293129085912, -2.24775674148539, -1.38839841727632, 
    0.395863905233043, 3.176755000392, 6.41394530815346, 9.32939998983173, 
    11.53752497863, 13.1878659063775, 14.0363587856162, 13.2063612998074, 
    10.2826431132315, 7.04445804397932, 5.49836289444132, 6.31700025929695, 
    8.28023882880633, 9.53125363412662, 9.46636280405579, 9.4139908776618, 
    9.87721338557378, 10.2531402484171, 9.63222516309714, 7.96099259968354, 
    6.29700607037049, 5.91162539375063, 7.10797565119502, 8.39497730694285, 
    7.96794256442177, 6.37501844733081, 4.64282778908115, 3.33556953195663, 
    3.02284149050042, 3.87712873738655, 5.70947134613352, 8.18119158407792, 
    10.3146679279898, 11.1508801884521, 10.8980568150134, 9.83313651969723, 
    7.64916163082465, 4.68999527349859, 2.2360186209877, 1.60369619024796, 
    3.29585864910954, 6.53567876985078, 10.2634584384539, 13.6924804608011, 
    15.999867203826, 16.7837933284536, 16.0898912284249, 14.4276707700985, 
    12.3689489780577, 10.7758558032455, 9.73320538662771, 9.21086997700739, 
    8.698245992014,
  10.3105245627848, 7.75412807148317, 5.96008645335427, 6.31699160049298, 
    5.2651848240198, 1.47119985097197, -0.892256663876421, 0.463959200059019, 
    2.43390502380925, 2.35248571455363, 1.96978059622682, 3.42778876715505, 
    6.29022569304271, 7.72557377052302, 5.51800893798675, 1.3925812567464, 
    -0.645451021500619, 1.04241604871834, 4.54272247657787, 8.26499489806116, 
    11.4838731245357, 12.7805002410096, 12.8577926232729, 13.3769655124434, 
    13.4843908999666, 10.7725633137203, 7.47129537705172, 8.245789882165, 
    9.40914325461888, 6.45162940994404, 2.88955666996083, 2.53643741138279, 
    4.21775069092039, 6.37055329759816, 7.92802123920615, 8.24597439524418, 
    8.32557388231078, 10.0775142677991, 11.3708930819256, 9.81884062648713, 
    7.29628545466934, 6.33329824530959, 5.48269977414056, 2.87888004856959, 
    0.790939219781317, 1.695924340273, 4.39538160488843, 5.8151466768591, 
    4.25911482632713, 1.2839948138016, 1.228852497735, 4.90060006346541, 
    9.50770027787785, 12.2632989896318, 12.6525884497942, 10.4357378745855, 
    7.13808439457296, 5.56345658087705, 7.08594518738077, 9.9321069518773,
  -0.142393924866818, -0.022257267507383, 0.266312682888241, 
    0.0156947646865673, -0.623010347454465, 0.749805112426262, 
    2.44124676921942, 0.147658305018708, -4.44361430716762, 
    -7.02369058659665, -7.93147465402821, -6.74302707627642, 
    -3.90706717455143, -2.68636965674582, -4.99078026894825, 
    -5.60371528121756, -3.29368755057726, -1.20123626828938, 
    1.02187650755297, 1.70201572734555, 0.997545822862932, 3.43093218574057, 
    5.04914083351114, 5.65565225994516, 6.70057114258497, 8.12900177628783, 
    7.66927284989054, 3.59044183103155, -2.40037647483291, -1.56042759560341, 
    7.9316245241352, 16.4311135039402, 19.2076223056194, 18.1956159831698, 
    16.946034387202, 13.1259500154329, 7.15273728953589, 4.03862323123184, 
    3.83608433085103, 3.82656961301646, 2.15967495780961, -1.3515115740794, 
    -4.60622941447461, -5.06631085117619, -2.65201742055376, 
    0.00354602389576786, 1.19586362317877, 0.784390340469183, 
    -0.504445958443494, 0.502359743660193, 4.11341107235121, 
    5.48598388260284, 4.4088202511239, 1.79065308256122, -1.3146092022013, 
    -0.532340383815348, 2.53043610304768, 6.44223101972032, 5.16011174225115, 
    0.913345975283631,
  -5.04207754125746, -2.04120957295356, -1.46444121163141, -2.11392877014422, 
    0.243656248037362, 2.84873028232751, 2.60339638729342, 2.21885569282409, 
    1.68289457723683, -0.800536327666131, -3.60774181833944, 
    -6.72347379196162, -9.88544530293049, -3.79519741256723, 
    1.59249418309939, -1.17475368766322, -1.29252772240621, 
    0.429818204811377, -1.61863369690184, -5.32112456306243, 
    -5.15727543690685, -4.92439483189292, -5.53683122592323, 
    -4.40551155533587, -3.55895160906971, -3.35676881864653, 
    -3.76587971304566, -4.97787649046866, -1.9057236552349, 4.43569185056868, 
    6.56012537903792, 8.44147614254119, 8.57227128058546, 3.35160259247573, 
    -1.43255628994462, -3.45189793482872, -3.86672560427095, 
    -3.89725364187238, -4.4501071952632, -3.14582726731554, 
    -0.908547748619928, -0.0700871785056805, 0.138688431410127, 
    1.11957613170953, 3.34650807386249, 5.70111792935754, 7.38620201846391, 
    9.903923333987, 12.4125660360105, 8.19797228820267, -2.69740833969003, 
    -9.14225635048238, -6.51668667828616, -4.39174298403499, 
    -8.35638276217533, -13.1386073225786, -15.820614957915, 
    -17.4615949444856, -14.4911904268336, -8.88084850168177,
  -2.60789566466588, 1.8815704258538, 5.92474992848538, 7.19793455128748, 
    7.87193490628192, 10.1670574662915, 11.633906718451, 10.1170205292251, 
    7.42661462408945, 6.92242289397399, 9.48990607963842, 10.8339887453932, 
    3.65754466392574, -8.34357378441931, -0.0701915138131069, 
    12.7180623747364, 6.97112925836407, -4.74036725670296, -12.0850483921613, 
    -12.1290872856534, -10.2866567806927, -5.87975207622859, 
    -1.5867053170406, -3.43566909402698, -6.33102716100025, 
    -5.28394920430102, -0.941839284408248, 4.23816534231332, 
    6.12806099186499, 0.234634810152409, -8.32597047001929, 
    -13.2731020418378, -11.1200023610069, -4.59334265134963, 
    0.465927485575771, 7.1034065518917, 10.7750205946374, 7.41228892958596, 
    0.672797926107098, -3.90255918716216, -3.02913968750902, 
    0.78310642555819, 4.16654930172891, 6.19983006388273, 4.9390421598099, 
    0.711208121877939, -3.03152850814044, -3.12024099905393, 
    1.55625165203209, 8.68196257914225, 11.4490659071072, 6.05897467572539, 
    -2.80468195737381, -0.284767482932599, 8.31561849737136, 
    9.53236922349246, 5.57697438251321, 1.39663965477446, -1.85000556180883, 
    -3.99523405521052,
  12.6512614611082, 16.3271107543132, 16.1247621025654, 12.7009402746058, 
    8.86557433139386, 7.54481700235768, 8.74188144623279, 13.6692112667381, 
    18.2244183837339, 16.7479664622461, 13.9336411709301, 13.9962341160296, 
    16.4935409243531, 13.4885410246471, 0.484537910661677, 5.48487372436256, 
    18.2861636423703, 14.2361609189432, 6.72027033672094, 1.17662520608143, 
    -3.49637249669386, -4.82671043267603, 0.301604132780388, 
    6.40783566829253, 6.23936411347568, 2.33271323023292, 1.5110818922068, 
    6.72044752707078, 13.718386186716, 19.8060904406422, 18.2224701058227, 
    7.0728729941187, -4.93834770234608, -6.91604763276928, -1.58736094429263, 
    3.87706040785499, 10.5602206560556, 16.1605814669562, 15.4987850016291, 
    10.2805545758198, 4.66696754239347, 3.97169781659544, 6.87334503291968, 
    6.6788240703165, 4.00427463581125, 1.38155150566326, 0.624007114431403, 
    0.917715834828531, 0.335930136848705, 4.31326310175386, 9.91981772321923, 
    10.7054760501308, 8.72884002073065, 3.02655382043305, 7.25775069584667, 
    19.3561259899376, 22.8944984643085, 19.235230604873, 11.999278086654, 
    8.5731918320265,
  15.7833437199672, 17.8961088253172, 21.9442638828204, 16.8312886211729, 
    11.6229525125175, 16.7794932146314, 16.2976162906395, 16.4051577654551, 
    18.970115450117, 15.9945419062343, 18.5611846297867, 21.361226480418, 
    17.5144270141291, 17.2476560609751, 18.3201458460735, 15.4989642893209, 
    14.1704353291979, 18.6763151796614, 20.9553645751027, 19.1015915808166, 
    21.569149202621, 23.6091229999786, 19.1483259885355, 12.2053180116805, 
    8.65754611763172, 3.76840555727567, 0.969746433508122, 10.5229373588276, 
    21.2548777448129, 23.4171854183919, 22.7325797906771, 18.7361008556141, 
    13.6860299668262, 14.6300266482268, 16.4955375647209, 16.4953255939552, 
    14.3832216538097, 14.5333956113547, 15.0026227225947, 11.8270256023602, 
    8.99055475089054, 9.49859827510205, 14.5649382555981, 21.0719452166887, 
    19.5118416577432, 14.3067362379482, 15.4864669103488, 19.9939963129531, 
    19.0689653971977, 12.9699835133985, 11.8342154181475, 11.288392403604, 
    6.52610503415561, 9.42873864892499, 12.843417737459, 17.7216560877622, 
    23.3442182231655, 19.5034763552489, 15.4238302764845, 16.0739991961186,
  24.0146466344556, 26.8309489696564, 27.0739571382551, 20.7261421500704, 
    19.3164684467949, 20.7550100992521, 25.896258079071, 26.8694831596968, 
    22.9024386387824, 24.3941988165799, 21.4990331596796, 20.4679298485563, 
    22.8995940978169, 23.8311086093311, 28.885796357586, 24.6359174842158, 
    22.1076750423983, 26.3450533332872, 22.0066534486095, 27.1910270562862, 
    38.2062912467798, 39.4708127814516, 32.6039246994303, 27.8583827931916, 
    23.2788416354925, 16.1125458222788, 21.1562452792407, 28.8410079472593, 
    34.610905223522, 37.1395516874487, 33.790400708428, 29.516008800175, 
    27.4409099763302, 24.0132790451693, 23.5691010673334, 26.9546002837381, 
    27.5840090892893, 25.1727847720294, 17.3696183207811, 13.0413939926645, 
    21.0034579170523, 27.5247175863577, 30.0701019853347, 29.0966094172896, 
    24.7135885793946, 21.800801856237, 22.7367101274095, 21.9058712942634, 
    20.9336048321525, 21.8013799942993, 20.9152183912826, 15.3250659895783, 
    13.4902561077437, 19.6161575322205, 25.1404809522408, 25.6072223927975, 
    25.7040582622665, 21.2391599537621, 14.2527847989143, 20.0623550069786,
  23.6448040224884, 25.1163030669365, 19.3547365134837, 16.6275558712242, 
    21.0202461777492, 20.2859061542434, 20.895847186134, 21.2040847074654, 
    19.496387184974, 14.4556661302868, 15.2595430886955, 19.101834756927, 
    24.4404123515481, 32.7512497210564, 26.3828950937756, 19.9499413018577, 
    20.601956226833, 11.6274325249876, 16.2039563538317, 25.8889345378624, 
    39.3915441365456, 48.4143231671183, 35.7016064829304, 24.508911297579, 
    16.03374678947, 19.4897713440333, 34.0458907535857, 34.5686441653588, 
    25.3493363549171, 24.4293726528318, 27.405400743208, 22.9912460127951, 
    16.6489197070665, 22.7904369203144, 29.0979704265409, 24.6959928694842, 
    26.2350558448646, 29.8322781966197, 22.7254205372897, 19.7498338706331, 
    21.7157870137086, 24.9322125447099, 28.3267943972117, 29.6226129154439, 
    23.5506121766649, 22.9049348861069, 31.1297177711266, 30.9582754035141, 
    27.5054080711328, 33.8197658315937, 32.5480610151666, 23.1431829663881, 
    26.0534903445363, 28.2526299292496, 26.5810787577101, 27.2785639768743, 
    19.6935922818345, 11.5377420114412, 15.8748256790079, 22.7713647872583,
  15.9372677851898, 8.9350926587893, 8.08414814542106, 10.3243763847224, 
    14.4905866247452, 10.309107671682, 7.27830316590666, 7.97707518892519, 
    7.27368831008451, 6.82467528997718, 14.0324111968123, 16.3907884626065, 
    12.7308721983141, 6.0202471657971, 12.0095769658083, 15.1918881620355, 
    -0.0966390771792312, 6.09001328766069, 27.4457827972527, 
    22.4260849874426, 5.232208130604, 5.08279754951681, 18.0144691738233, 
    13.2974629391941, 7.08214019229839, 23.4309147749331, 26.0376322811141, 
    13.0903509791224, 3.68441685957417, -0.846785244686707, 
    -3.19757815735673, 1.82212193734885, 18.7600839788871, 25.3463145663736, 
    17.4389413655108, 10.7373322431313, 5.87983940455603, 3.99232184638047, 
    9.39590253560308, 10.9332229128889, 14.1409350787184, 15.7227901288107, 
    4.3952913258006, -2.36088127335598, 5.13698230865648, 19.8993383396642, 
    19.2175646122822, 14.8450394659294, 11.3668630215254, 9.97232463420635, 
    6.48050495388123, 6.42274370339758, 15.0765522477081, 14.9409705487193, 
    5.22985035079622, 0.901200520160808, 3.37131775983711, 14.106398534554, 
    23.5937431179854, 19.1349558216827,
  0.276571489797525, -0.697721679230103, -2.55782586888867, 
    0.297824498779838, 9.8630509766386, 6.39005001457198, 12.1717929582295, 
    4.29074750370063, 13.0361303747982, 11.1640699331158, -1.23396521900452, 
    -1.97113247100274, 0.90425303046605, -1.03264473072538, 
    -9.44147568200494, -9.51275120869717, 13.7786952610387, 26.8200487400898, 
    2.54375830855036, -12.4355450324782, -8.56797259722366, 
    -13.7610510211859, -11.617957173378, -6.6677953634133, 15.3343068209976, 
    12.0698266418646, 1.77835678516522, -6.36092871015797, -8.19633432924467, 
    -6.30067448692788, -1.09008711869874, 6.70425200989285, 1.75036344277887, 
    -3.4886275950862, 0.241499746159465, -4.14801633468354, 
    -3.67534323009684, -0.849538938992662, 14.0772668991345, 
    23.2449519081357, 13.3558089955788, -0.731119578672761, 
    -0.845277943865706, 6.05224451472602, 10.7739992556753, 
    0.691663899289959, -4.67548655608955, 2.66649122432173, 3.9275988260674, 
    0.0878734548839608, 3.51906606528062, 12.0487372012505, 6.16625537040846, 
    -0.94188751520991, 0.166306206937946, -0.272756737067445, 
    4.49812708222489, 12.3881354252651, 9.7499070802299, 2.16390931292587,
  3.18916638006775, 4.7810770542431, 9.85405907290891, 7.52695665082449, 
    12.5165122982429, 13.9020287065915, -10.4578992985522, -17.7782478976273, 
    -7.69253623430893, -0.545593104984474, 2.90484769700138, 
    -0.87687950737239, -5.8998704667362, -9.26130349117428, 
    -1.18592557303792, 15.855042603856, 4.40748857254822, -1.7551809673252, 
    1.02768664417901, 3.36346564506848, -5.70568338659752, -24.1343459939312, 
    -11.9754758711666, 0.994956255982859, 12.3947595744414, 10.1503541603356, 
    -1.20828953020111, -2.19083387690702, 3.34148415187587, 7.33946743004682, 
    6.15973281344695, 4.0666366265194, 4.16901670513572, 2.1310748153896, 
    4.39625865371857, 6.8263617639891, 8.27095633704817, 6.18628338644648, 
    3.32765001672415, -0.0498234559393965, 2.22695160510386, 
    3.46835345516811, 3.14090918293011, 7.5130436253434, 8.26645172372194, 
    7.55294994045049, 3.87487673271667, 2.13091893218329, -0.233464784632972, 
    -5.99461182795536, -1.86681746299399, 3.13430411240914, 7.42522322585048, 
    2.57071900638021, -0.432003473492072, 1.46677457219229, 4.90942840826959, 
    0.0293796002701661, 0.253016614386317, 1.58695560918747,
  -1.71898511055433, 1.66999484381081, 1.53793997831149, 2.97601044071168, 
    1.30186564432685, 0.152227689937618, 5.90964542330908, 8.98469218111136, 
    -6.06647444288842, -8.39816362064031, -1.5430117933868, 
    0.173611728221627, 0.0171056953323042, -3.10604713113046, 
    -0.707386707724115, 4.93802058040027, 11.0973617752464, 1.56216014581256, 
    -0.513149739737826, 1.10389946018384, 1.4779867502612, 
    -0.974540716258676, 2.92786222346692, 6.63324375994838, 9.13662535373996, 
    0.980394495781619, -2.09501437913958, -0.937771928116349, 
    -2.43298622578366, -3.2885226774732, 0.530064745717073, 
    -1.24762512598094, -3.96186922776581, 0.62052820440237, 7.1020139823927, 
    9.55142303690895, 7.47031028732721, 4.98532888423554, 2.20932415747561, 
    1.6182082536214, 4.60513639142845, 8.06739055916096, 8.22360763415698, 
    0.289678270316957, -1.42275595230699, -0.16440967134321, 
    -0.0362102405999289, -2.22501370563064, -0.338881483570395, 
    4.08372718094555, -3.77636329511697, -0.464957282934408, 
    4.03906473309219, 4.96311759272753, 4.8823802070683, 1.5860519213327, 
    2.84690867323405, -0.0826580584435572, -2.60526149959429, 6.35713044210165,
  0.0318995282050722, 2.95971582318827, 1.72737519886796, 9.67161230874551, 
    11.1939332393139, 5.03943952851218, 0.620838142457469, -5.81282857513502, 
    4.96288672512594, 0.2344858756717, -1.23438806391043, 3.43849805732832, 
    9.24533636263191, 10.174603634836, 7.07848169164803, 4.98379028187784, 
    2.53510202726085, 2.63558863278038, 1.39259232958259, 3.04046836684895, 
    0.990816905576068, 13.4287765146216, 16.7275734039729, 8.2235776026296, 
    7.32169157575164, 3.77015488417904, 7.72107608059147, 3.34784317889618, 
    -0.204734123998291, 0.76788040095151, -3.77029304453594, 
    0.532054070908363, -0.799139218903216, 1.59519433886022, 
    4.53719641499754, 3.86012596410818, 4.37063093740194, 7.35799207964609, 
    6.34043933283871, 3.91423856973872, 5.84547722011939, 7.06231289728193, 
    2.28840738239162, 2.65852106456765, 3.17606133974327, 6.13561482447806, 
    8.36014247075756, 4.08866314834728, 1.71897946103789, 5.92425144042928, 
    6.11044617359288, 7.03235267998186, 8.73457365361088, 6.06052430250552, 
    1.15798304988936, 4.86327164895006, 8.31096450701644, 8.12815891233472, 
    0.20248012366748, 10.2971991991183,
  -10.2812326901392, 4.0671897940107, 2.67463415529422, 4.79346873589, 
    8.32495152590625, 8.11409813908086, 5.84200924414545, 3.71922966609402, 
    9.81387358782872, 14.4698580147229, 11.477249184317, 9.10660798608432, 
    8.78018299419643, 12.6850209317342, 10.4706028918568, 7.4942685914536, 
    7.2563337314677, 8.66204023852131, 12.6596972891751, 11.5020403124131, 
    5.53994022252859, 5.40352238726006, 8.98849543188168, 15.3734449688462, 
    9.61803705836262, -0.288018901665395, 0.366633354464334, 
    8.16211826654979, 11.2628741462068, 6.27970925573561, 11.0759793176953, 
    19.1010713047145, 11.6190264467014, 2.76911219506262, 1.92031970032256, 
    -0.360534654615619, -1.82572584634991, 3.831647295508, 13.158254390054, 
    15.2963652262741, 12.5432613990738, 12.5410012409807, 9.66911783770297, 
    7.51774585057743, 4.4848632307734, 5.71053537969165, 8.0751593623602, 
    10.0162823528439, 8.54354265949395, 6.33232368010832, 8.87503274673476, 
    10.943361751104, 10.2720817898736, 12.9606454410174, 14.0543600792915, 
    10.7452513455826, 4.48303805692279, 4.91767563636965, 8.27342793071171, 
    -5.44889304799508,
  5.07873429123313, -2.88722490435298, 1.88720926345098, 4.40000231190142, 
    -0.674447004773608, -0.25231274030432, 1.84380452590376, 4.4626151147038, 
    13.4017691009862, 19.5333718305775, 16.7502868508744, 7.96471815427271, 
    0.292983661398295, 2.09293206904913, 11.3554377568949, 13.0203318334, 
    6.35922199827673, 4.42326110953396, 8.57743630013047, 13.0820007114996, 
    13.0231588403541, 5.74340487544547, 2.12991956928146, 7.18705962852846, 
    12.2810852275898, 15.5446009461816, 11.4706844469261, 9.07803631677756, 
    12.5877669645742, 20.4404389027263, 15.9387200035685, 12.2584086579906, 
    17.0765320571911, 6.60319960290683, -4.29821880089971, -6.60826781859864, 
    -7.95166014735433, -3.75594018209222, 6.67143022804934, 17.6614374369705, 
    18.028172436887, 9.12543536205943, 2.35907066349816, 5.6183623831311, 
    8.86869882983012, 9.2897773902538, 12.0187542462603, 14.0513360544119, 
    10.6311537080056, 12.9400598786841, 8.11835810784516, -1.79910900566736, 
    -3.54929390337042, -4.75584016565376, -4.76651140745249, 
    0.213340128464938, 19.9299646915726, 22.3930233497513, 20.0486241197149, 
    15.0585029160748,
  26.8088279729391, 29.4539925013601, 23.1538591272227, 23.2650711800095, 
    20.300134044752, 13.229189608807, 8.94206543294252, 4.2489907739086, 
    3.47245839256703, 10.7690143323961, 20.9491968216598, 24.2634161988362, 
    16.1599130025903, 3.3475891941735, 1.06406177753737, 11.9447879509948, 
    23.3773638388342, 24.7321840539295, 15.7634067052926, 6.75403123456838, 
    6.80859454147987, 17.6698602436099, 20.2393730545899, 14.0751078713981, 
    6.28785604915141, 7.93286373456791, 18.2607262690883, 22.3972270012233, 
    19.9497562991592, 18.6237822528367, 19.682073341615, 17.9533704517385, 
    19.0745873018314, 26.508216369962, 19.4710701212964, 9.6300481540474, 
    8.95792876479511, 11.163278568485, 12.3886724208492, 13.5009326382389, 
    17.4220037331179, 21.2836894499426, 18.9417107955864, 13.9412974219063, 
    11.5158202736256, 7.83226644713247, 4.0225389240073, 11.6275156342839, 
    21.8448645093571, 20.8942954227443, 19.9512628951983, 23.1860063285201, 
    17.8966823623303, 12.2341248827733, 12.0364787313609, 14.8436463438657, 
    14.1639724607924, 15.9756832178936, 28.4354274882206, 24.5197325030285,
  31.8220738785871, 32.2052324301498, 26.3261152791381, 20.256606728553, 
    20.6483044485339, 17.81198013201, 17.5939197073574, 25.6805251253144, 
    27.93747167006, 20.5570445420568, 22.0040426220269, 26.2742343968312, 
    22.5418780357412, 16.8045571028726, 13.154084958604, 14.6717153560537, 
    20.993508830116, 26.7867004459784, 22.0639228376356, 16.9688381124511, 
    17.741044824739, 15.570482165049, 15.873450923151, 23.1109587621117, 
    29.8907324763338, 26.8030390798898, 18.3825551317621, 17.5396119120873, 
    19.9134191515809, 18.7694990144869, 17.3169336006557, 17.2802904801147, 
    18.7116256076612, 27.2317419420365, 33.4043385288485, 32.9299244238867, 
    29.8469546311212, 25.1052168042731, 20.9464860304787, 18.6854289996882, 
    19.3563394814181, 24.8681043892724, 28.5351682150129, 27.307388349216, 
    21.1308339068065, 21.292334128032, 24.393333053209, 18.0082306981931, 
    16.8203686210261, 24.9450232959165, 25.2066614054399, 24.1881184546466, 
    30.3641380935251, 30.6183738049036, 30.3712147453413, 30.6554346120855, 
    30.6179594691557, 25.8666177421415, 24.5180777148846, 29.6153659826476,
  18.8332715118931, 23.274863235146, 24.264351906627, 25.2517805943889, 
    29.0204446046619, 35.4984552358749, 37.8709458734988, 29.0512642102521, 
    19.6520369817795, 13.5026109059649, 10.9916143937192, 13.7984779865973, 
    17.6167497457682, 20.9818510795681, 22.6159776084258, 20.633288988712, 
    16.477230185286, 17.951349112244, 22.1640826415808, 23.3566465746787, 
    23.2419136873267, 25.2944979743028, 21.8494433447937, 17.6129241391931, 
    25.1539274462485, 26.6158770284814, 19.2574106238738, 15.6289526290818, 
    12.963464636433, 14.6497403220539, 19.8328161777465, 21.5295183566299, 
    19.192367698501, 21.5799104630555, 28.6555532892007, 27.2738085375254, 
    23.2234247202182, 22.2727158123409, 17.5920985024393, 13.0492813615134, 
    13.6731992002421, 16.5073378297662, 18.5477938521792, 19.8732307811705, 
    19.6568733995615, 17.0469712975764, 16.5638000923247, 17.2450882559416, 
    17.2226464299129, 22.6345177469929, 26.8214080211052, 27.2917732601751, 
    27.6516608585287, 27.5613694348308, 25.94091983614, 20.9273771527616, 
    8.06718153616945, -1.91048273224047, -1.92646984415273, 7.95137216905338,
  22.1329950813489, 21.0264481066714, 15.6791704509726, 12.3597654051879, 
    12.7922476542236, 12.8449727018773, 11.4188853250537, 15.6902236552903, 
    17.9766924629288, 11.2416675583279, 3.37615344388047, 5.47640081462142, 
    11.6625419340388, 17.0465021901277, 19.8095882672988, 13.2418886038269, 
    4.35376338373179, 2.66005720775822, 9.01634860908546, 13.0294711207901, 
    16.2152415169821, 20.0850480867593, 18.2969466587704, 17.3047399435542, 
    12.1812463177537, 6.56165884604687, 7.69234905429868, 5.79875839641672, 
    5.77673142912899, 9.15363319271606, 9.29689822775303, 8.03843417332958, 
    5.13504509779771, 3.00956789117056, 4.1566918464592, 9.06651988140799, 
    17.0825221124065, 21.3932447611458, 16.2184533379215, 8.0971625654004, 
    3.45694696140451, 4.93646024702824, 10.2666924754015, 11.0351552855842, 
    11.0642608690164, 12.4080397352249, 11.6575380563442, 13.7012181251496, 
    18.0537206756937, 20.4537802197522, 21.0776453006316, 20.866824669126, 
    23.4298505996556, 26.2977382858782, 16.2667226450459, 4.40998101746424, 
    3.57092529099666, 7.02146388227865, 11.3662711408925, 17.3308737326965,
  -9.12757766867846, -11.2855173695976, -8.27667731002669, -7.71783592684231, 
    -7.45220113805092, -1.11514368178124, 12.104057671366, 16.3711626103413, 
    7.32545414414035, -0.590641468118274, -2.17060731608505, 
    0.449224278781446, 5.64632982196027, 8.94063831178632, 10.0075217112716, 
    11.3587546477969, 11.7876282198511, 10.4923616666273, 7.94234628789973, 
    11.574192950108, 22.0647003138019, 21.0691532898302, 5.12325289713992, 
    -7.5433590138906, -6.5789064436835, 2.98888827160259, 7.58463194655241, 
    7.87040675841733, 8.59418004482815, 5.73188974290618, 0.317355002240704, 
    -3.25723885139893, -4.94156942885038, -5.03649993994964, 
    -0.394933886656375, 8.97301917180122, 15.5451884159535, 14.1214539334529, 
    9.63671268460229, 6.80027756990366, 6.56865925221663, 3.61630769557229, 
    -1.81967084067115, -0.0305374255194656, 7.38070051764775, 
    11.3527432403129, 11.8293481138113, 8.07012063249401, -1.33740831994585, 
    -7.25598236763875, -6.71134502922619, -6.31922279649346, 
    -6.99823687617974, -7.24838662035442, -2.32096489731627, 
    4.89120367938282, 7.66399388932005, 5.5107229249462, 1.80996070307841, 
    -2.75332398724245,
  -0.0632815697346074, -3.53885720314941, -3.84668206058873, 
    -2.2177688840255, -0.0229042636461103, 2.81008639216484, 
    1.30093817126593, -2.2214647849869, -3.13260413780066, -3.16436701676677, 
    -2.39115051799796, -0.175008197339484, 2.20705994848664, 
    4.57827378909538, 7.35928471445054, 8.8241628492779, 8.79481271862646, 
    8.21219293235625, 7.38617096986089, 4.06184910290174, -4.32348127591856, 
    -10.1317519645193, -6.99925943720577, -2.05765328435429, 
    0.40280683670224, 1.4680061909323, 2.92622442649679, 5.72412101013594, 
    5.73463841210012, 4.1708873258608, 2.82491983964019, -1.5084382224781, 
    -5.95202408384474, -4.46282984561038, 0.719590252321036, 4.0813338837487, 
    6.5122705431311, 8.90831593983518, 9.335789215861, 6.29518968707902, 
    0.482099251222314, -3.53326452677032, -1.78965217383736, 
    3.28543861433127, 5.6367433879887, 2.57428257011561, -6.28663463960225, 
    -16.0196703094613, -16.6626001181238, -10.2341907384683, 
    -5.41135815800596, -6.05255686705668, -6.15913249881718, 
    -0.606624710090902, 6.28955796979436, 9.3043754574873, 8.38048964518213, 
    5.0619890450936, 3.01718732989214, 2.30283823593556,
  0.406912548503223, 2.95474411661435, 2.29124739745102, 0.0787802225187181, 
    -0.4985092300662, -0.131583001558587, 1.15231602349655, 2.64907520323633, 
    2.83726209730878, 2.21637651550535, 1.25089795763809, 1.58007755751712, 
    2.18903541352581, 1.30154961276641, -0.251515536489114, 
    -1.60445238678262, -2.32143066399852, -2.21504796116716, 
    -2.04077299859735, -3.4006155100576, -5.04199497413399, 
    -4.63728175460375, -2.92144583367355, -2.47875049340359, 
    -2.63316318882658, -2.09388342616575, -0.655523878551981, 
    0.824114606856427, 2.16167511917989, 3.91729491891702, 5.78533014232479, 
    8.75662958368213, 12.5979303599742, 12.5036970274356, 8.00771508406717, 
    4.24201503936332, 0.300817675724487, -4.63494125183102, 
    -7.02234789454254, -8.48351822587656, -9.4101504413407, 
    -9.84594200720944, -9.14027506219829, -9.82614347437498, 
    -10.4367764374031, -6.54941052894183, -0.235573158342821, 
    5.60223927722813, 6.45953232240895, 0.750227719379027, -4.82871766573973, 
    -0.760549393437916, 4.77452716514599, 5.30336403067089, 4.05839948193201, 
    4.31632389610087, 7.26579762567421, 9.25031544014492, 5.63399134405262, 
    0.469333602227834,
  8.12811781006167, 7.87647347249121, 6.71997852235946, 5.61496740865235, 
    5.44222330175093, 5.3517433446565, 4.00054603097583, 3.55227532869866, 
    6.12115345123199, 9.71221926963587, 10.8264264145372, 8.98947999442744, 
    6.09018638311639, 3.60339051990647, 1.42097291655491, -1.45234629756791, 
    -4.62594815542258, -6.55052861438321, -6.34370075019669, 
    -4.31794546381421, -1.85710538893769, -0.277047981455016, 
    -0.375720259023724, -2.05485328932117, -4.22452511086121, 
    -5.55733413576393, -5.53188374856848, -4.19858344618176, 
    -1.98169248765748, 0.540810880125252, 3.55394053531595, 6.51600145294947, 
    7.82930924410164, 7.06022870000503, 6.16933250863292, 5.60163270536153, 
    3.61841430283247, 0.891703204481862, 0.0419178700671357, 
    1.30600319821428, 3.03800865709758, 4.46936719169542, 4.57348061653108, 
    3.18099640994672, 0.965123084622324, -1.77119807343904, 
    -3.20834989454139, -1.22188630022804, 3.4154407593857, 6.83242910435291, 
    6.32067934731511, 2.39940702676052, -0.555194537507283, 
    -0.647193089691669, 0.865861444276197, 2.86076830098839, 
    4.46023879129661, 5.63175163315912, 6.43298935820573, 7.35339896864189,
  6.31145542946035, 9.50785574307717, 11.6812237842749, 12.5401600258304, 
    11.8804896943129, 9.72694163759745, 6.90072625958547, 4.86300528136036, 
    4.55040121321974, 5.99354424343129, 8.46691421087225, 11.0191532858538, 
    12.9797164416586, 13.6865401496439, 12.6167493163444, 10.0273470008777, 
    7.3509733013912, 5.91987261214991, 5.33130497881241, 4.71145941993891, 
    3.67057293724687, 2.61831453592438, 2.39481047543397, 3.68479563336175, 
    5.93739151582831, 7.70945951222793, 7.75853370030457, 6.15222709476731, 
    4.32958235876149, 3.53415414959401, 3.57137836795393, 3.61978600523052, 
    3.30142673886842, 3.16635405442697, 3.24126129783155, 2.4960747505967, 
    0.659670487319176, -0.571130155277361, 0.956661123879681, 
    5.64627130218721, 11.1762234213553, 16.0625058242951, 19.6186716401869, 
    21.6200172454726, 21.6266484981363, 19.570572837214, 16.3307121875537, 
    13.2019332072747, 10.9552871288107, 9.84970905311868, 8.39811335285531, 
    5.60225603582237, 2.45778410987094, 0.340716582818907, 
    -0.588130195979869, -1.13923880655812, -1.63409477309266, 
    -1.44182116878521, 0.0246609672158114, 2.76796155195319,
  1.70819520886991, 2.17207838640878, 3.59712739898449, 5.36841338993652, 
    6.69450144137824, 7.02992798187749, 6.32283282597769, 4.88663437827509, 
    3.22957116948168, 1.96073502791653, 1.5100057809024, 1.79957345647494, 
    2.34483759259596, 2.72328249755111, 2.79068310873644, 2.88137280129257, 
    3.49366051944615, 4.98109061467992, 7.29882348216543, 9.87330544884735, 
    12.1903925755801, 13.9367054647857, 15.0874421381073, 15.759729388819, 
    16.0241917048683, 15.7726274004165, 14.9009468017632, 13.2183228887161, 
    10.8001777424435, 7.96770250997837, 5.34118108236705, 3.62459842294564, 
    3.27554945070887, 4.19162941339372, 5.86237461330023, 7.51228158724563, 
    8.54684355198768, 8.94906007472621, 8.88832403779088, 8.5523867188657, 
    8.58050599912972, 9.16348929619478, 9.8979654420353, 10.2698684583643, 
    9.898846660319, 8.87175149567225, 7.66056664607468, 6.79266928469594, 
    6.46281209712639, 6.69623463811391, 7.33013898632247, 8.29804752350733, 
    9.35184169115979, 10.114257913551, 10.2042661813585, 9.33730057542303, 
    7.79173499110352, 5.99762910376274, 4.07871137070369, 2.43700932902005,
  0.69530563339694, 0.245758860317243, -0.0852140000111819, 
    -0.298560786384749, -0.410162151736902, -0.443936133007234, 
    -0.418099402152881, -0.337383908615291, -0.195025466718228, 
    -0.0439777626138378, 0.0563842673241305, 0.118827955295367, 
    0.209175543724457, 0.364592415970481, 0.617245522029146, 
    0.998322781357695, 1.48447048042215, 2.04312410030206, 2.69122372432333, 
    3.43623720771197, 4.21635139563982, 4.97399401223729, 5.590055933727, 
    5.98946366873222, 6.08140446257038, 5.82347620257587, 5.26404452917703, 
    4.47112669919664, 3.43933677059567, 2.27341484629534, 1.17643973819881, 
    0.32951962937464, -0.227486491081089, -0.492385014496216, 
    -0.504124343562125, -0.323665173980832, -0.0349720147092489, 
    0.303637082299958, 0.616403826805444, 0.826838511018993, 
    0.893560984158534, 0.821160868108026, 0.692268923371942, 
    0.585147177347042, 0.54570077474896, 0.615282972265947, 
    0.784797446674624, 1.02390589744034, 1.28051284521228, 1.53416019033826, 
    1.83012355795717, 2.13525895567941, 2.38678411813175, 2.55474108117634, 
    2.58813124260122, 2.45136344241914, 2.2422540043386, 2.02277093076492, 
    1.68925962411165, 1.20731832455686,
  -7.15178415153569, -6.91162659288842, -6.4658685995786, -5.79500151017961, 
    -4.91870268244903, -3.85463206180315, -2.69362359915054, 
    -1.54760568206488, -0.494555553775476, 0.438490579621445, 
    1.2273894293286, 1.87383421258163, 2.36063297752798, 2.7064204573759, 
    2.92510396151275, 3.06070771287394, 3.10300444452984, 3.04793238814465, 
    2.90664371938474, 2.74704131504129, 2.59276816610013, 2.36807310555286, 
    2.09957746051724, 1.81903110115797, 1.59039543910108, 1.38352368091702, 
    1.15180005933456, 0.88243455761893, 0.50750762345025, 0.0489682646338712, 
    -0.419353018482442, -0.896654032787862, -1.35060493705213, 
    -1.71700236478922, -1.95844836254201, -2.09596724577079, 
    -2.13144809226836, -2.06666676475696, -1.90525581610918, 
    -1.65371336719802, -1.30726382643723, -0.901689779159614, 
    -0.541662542990874, -0.270427066558619, -0.0334181686218194, 
    0.163186238880337, 0.235285567361533, 0.133483309869935, 
    -0.146687003726741, -0.598781859416999, -1.21646904429485, 
    -1.96847414937253, -2.8047187303743, -3.68206180965643, 
    -4.54022699832374, -5.34738900284858, -6.04903967439551, 
    -6.59671168686993, -6.9759372319528, -7.17125438124782,
  10.0842594966006, 11.2127370414636, 11.7964609666874, 11.5293319988379, 
    10.4476409916605, 8.83399296363373, 7.14979338469542, 5.69222802388875, 
    4.49534383682899, 3.5376131019344, 2.96546922916245, 2.7444888622598, 
    2.77067001052863, 2.91956388944311, 3.0934415459657, 3.2540642734273, 
    3.33917078375448, 3.41258889959601, 3.29621654016381, 3.34510315595889, 
    3.72224245029359, 4.0368018253746, 4.06405833526447, 3.67842124098704, 
    2.86169806419007, 1.78267194884286, 0.702096269771862, -0.16914364755983, 
    -0.573015694687622, -0.475683652500089, -0.0897500802626791, 
    0.315138552789754, 0.454539933260459, 0.158660161838202, 
    -0.552593368252541, -1.41655626490925, -2.05273261471679, 
    -2.12960476807183, -1.37055655503016, 0.186235081623633, 
    2.20477281732991, 4.20285633245331, 5.74419811711195, 6.43646803993577, 
    6.2463537750137, 5.46520788197797, 4.27177888909102, 2.84012693156535, 
    1.51368975673148, 0.586269994187505, 0.258473802391734, 0.53117853551253, 
    1.28048590776883, 2.41653912263599, 3.70156352552237, 4.86750361356895, 
    5.84749524557976, 6.70986949481458, 7.64048329732519, 8.78778801622273,
  3.96713984815642, 2.05661231587469, -0.254444600324911, -1.63277743095133, 
    -1.6572310644905, -1.13906137586815, -1.4039200355296, -2.1959846579831, 
    -2.44629807811411, -1.41486768178372, 0.486652316998422, 
    2.54341010958645, 4.38315000130457, 5.4518174558782, 5.8805305146371, 
    5.22406630935486, 3.43900716884821, 1.18777644272515, -0.822765343960309, 
    -1.44336316284849, -0.733760780695123, -0.383865815105977, 
    -0.215090985334183, 0.425753568956471, 1.53663047994833, 
    2.27430363798935, 2.13034615644517, 1.62782835123674, 1.47344400500395, 
    2.16136797499139, 3.92157415344098, 5.4635711128515, 5.53650234475684, 
    4.2990673661409, 2.96213434907238, 2.70645331926987, 3.82636010423903, 
    5.29415843509271, 6.40400910588948, 6.93821563086155, 6.87644346058655, 
    6.3417000374244, 5.5692297939311, 4.53355132051625, 3.11934524464782, 
    1.95336575957239, 1.74587488908176, 2.68189226046911, 4.41648746924217, 
    6.29272975295428, 7.90768435574168, 9.05624230788171, 9.05404440529823, 
    8.20775290971814, 6.89406358848029, 5.77616896738982, 5.24056870751065, 
    5.04240197414277, 4.98883361275554, 4.83138446300821,
  4.95833571143053, 3.04512053209861, 1.5242692433812, 1.65343943803785, 
    1.15353029605718, -1.32558758256589, -3.88989552200002, 
    -4.52576280442162, -4.39175331996643, -4.42773003049973, 
    -3.50150232520218, -0.555497406904755, 2.10822933378889, 
    2.18085743530524, 1.35439468753346, -1.49464629885566, -4.7200268054694, 
    -3.9609949670403, -0.455987144623191, 3.48184311901141, 7.07757023129652, 
    9.01302587325361, 8.97697373547797, 8.14142501275741, 7.0132132227662, 
    4.86071364738403, 2.34535137863369, 2.87802716406407, 6.03104974006643, 
    6.11697412678784, 2.0465768188482, -1.18017744958315, -0.679103765244666, 
    2.21965549329747, 4.88379886511139, 6.44908126334315, 6.77898823573407, 
    5.60192952380431, 4.13946831291237, 3.8812818872582, 4.33535246828487, 
    4.58735021021108, 4.16339523202686, 2.72515655489116, 0.75674419607936, 
    -0.111186213442482, 0.437393446028312, 0.491810642292215, 
    -1.59962745620851, -4.56953348659035, -5.05752802962012, 
    -1.25372748627014, 3.54574535540035, 6.75991781397021, 7.35335462986024, 
    5.49348949144697, 3.96702234870514, 3.22664225331946, 3.35712520782436, 
    4.66501489527346,
  0.216439105184341, 1.11057382719744, 1.74157705366104, 1.05743106361565, 
    -0.649938749460852, -0.738551030516875, 0.56163637402062, 
    -1.67837498687062, -5.83473303610957, -7.22956083277924, 
    -7.82181917492695, -7.9179774206077, -6.00865589864969, 
    -4.98901530621088, -5.80747626978676, -5.82676702076737, 
    -3.97260614224357, -1.4172024291757, 0.640632424261527, 
    -0.246363660213689, -0.0551528641063886, 3.41880530062089, 
    6.07456644962153, 5.12793971991021, 4.55983032400332, 4.07396762148926, 
    4.74389430332364, 3.69561133403456, -1.32127593870953, -4.46907960114015, 
    -0.446034583490916, 6.02498206956024, 7.74279775207444, 7.15228837340743, 
    7.02643498648534, 5.33244716227972, 1.37231353779934, 0.293179832272875, 
    2.51916732477397, 3.32393720373038, 1.65430165706007, -0.997725286371809, 
    -4.05998233626575, -5.50984700947076, -4.69208734350767, -3.251648983967, 
    -2.11279757950034, -1.45487028193671, -0.681192917324532, 
    1.55179144174045, 4.28238595262158, 5.93672131821111, 4.19114052760628, 
    1.41363941176062, 0.276398827381726, -1.03539470762919, 
    -0.337984996498856, 2.87236091911256, 4.04507890439899, 1.4129079023124,
  -7.48573249182509, -4.85239945264829, -4.31495787643369, -5.20625071021014, 
    -4.10777669854352, -1.79340465219292, 0.309621673064512, 
    2.59760280674227, 2.57531485683871, -0.885501534238706, 
    -4.35810362857387, -6.31975769387925, -8.20341582732698, 
    -5.50725152880154, -2.81120980198048, -3.80195927868343, 
    -2.22466575512694, -2.09562282937093, -6.50760130124151, 
    -9.57764285700196, -8.7399848583655, -7.84389356966631, 
    -5.94375025253555, -2.15981843731585, 0.0881974372258509, 
    0.404079182546137, -0.542552159548025, -3.88647754258912, 
    -4.9571243946157, -1.88394456661047, 0.0852382608785315, 
    1.66882511718676, 3.68564627344804, 1.85983921035962, -2.3137408120758, 
    -4.84248336581505, -4.51587064142081, -4.52565706401211, 
    -6.2174119968781, -5.78504737803167, -4.18342872525126, 
    -3.86412168089351, -3.64074273302645, -2.94940530080728, 
    -1.81148431112453, -0.847960470435904, -0.297583371160862, 
    1.22814795833027, 3.67283298692774, 2.78022132946633, -3.88429545593958, 
    -9.56593250044057, -7.29032048390585, -5.20357449701266, 
    -7.80612288415425, -10.1996063012341, -12.5366938434073, 
    -16.0466093255738, -15.3354601352595, -10.8171269169042,
  -9.56085960439344, -6.109494302597, -0.776974042204894, 2.06548859057768, 
    3.42621744705988, 4.78144383813922, 5.57409200205025, 5.85199244804636, 
    7.08351448061234, 8.82707131859022, 9.06224768319748, 8.32182367818094, 
    3.16338458305829, -7.02276908689884, -3.14504575504907, 5.34122359879377, 
    2.49403186939516, -3.91970750485873, -9.45916259141378, 
    -12.1473370477233, -13.4319514617428, -11.9820552188059, 
    -7.8045329578924, -6.955106380122, -7.14237453616734, -5.43470090505964, 
    -3.78379973631235, -2.09321613930986, -0.872458454654529, 
    -2.98010463647688, -6.68945778833768, -10.9469197609128, 
    -12.1010123903177, -8.59493248779064, -5.03799036892079, 
    -0.136781044903587, 3.43725001099737, 2.85155024052745, 
    -0.35781268065036, -5.17174926293759, -7.21116857763116, 
    -5.23477190356036, -2.65752518408829, -1.36750799789339, 
    -2.57473469130235, -5.31001124821153, -7.33372245908883, 
    -6.78105921297141, -2.41271302775075, 3.01133532328724, 5.5732296105006, 
    1.82862053935904, -6.74329824004398, -4.73863457427501, 2.85858089489669, 
    4.66432278540696, 4.691843783967, 3.90415173799322, -0.265788950768696, 
    -6.85162093410982,
  10.741623783628, 11.4671555107657, 9.4960527002808, 7.70492155932814, 
    4.23661166640506, 1.31191520568839, 1.65487830918768, 6.20996301289681, 
    11.7298074168893, 13.5363006116847, 12.7940603451459, 10.6589735323213, 
    11.5244156939363, 9.50704353742821, -2.28841104112311, 
    -0.0933844503117777, 9.7084443884671, 10.0461318626225, 8.55412360546929, 
    5.15439288608706, -0.710504996948722, -5.03490304673505, 
    -5.10801805937799, -2.27769851021966, -2.43139581292507, 
    -5.62274004137061, -5.98632614420361, -1.67803349511425, 
    5.50764622379669, 11.0708329514022, 9.63551363182383, 0.77463977188126, 
    -9.01398429885503, -11.6516121635993, -7.56133945552732, 
    -2.8825836876825, 3.65178362689029, 7.92876152657887, 7.82838341607795, 
    6.16040688138726, 2.43159000755952, -0.108508516919207, 
    0.456790751085519, 0.927563824200472, 1.05842383996767, 
    0.475887107297917, -0.195466823960273, -1.02477662259615, 
    -1.62086025679949, 1.81241021836548, 5.85291818760773, 6.73187340457635, 
    3.48115819082924, -6.06992650336139, -4.66583199654149, 8.07386447117004, 
    13.2856131398931, 11.4126682208605, 6.76676345847008, 6.33765809323601,
  5.83948247093262, 8.43322809319532, 11.9337555042912, 8.50914420408716, 
    7.05826210834146, 11.3904943717562, 10.9734992528151, 10.0813367072879, 
    11.2337918124357, 9.78652297915108, 12.889348021963, 15.9064083408052, 
    12.0355437005841, 11.1431256946481, 12.668407563878, 8.21430682315769, 
    6.81153541483791, 13.2460665132777, 15.984303226317, 15.7376457280839, 
    19.1562717497588, 20.3031960811486, 12.8814847459369, 5.67239451159461, 
    3.88879870568136, 1.05386188125136, -2.53741608176615, 1.61508947623233, 
    6.89044166849024, 8.85529400033105, 13.1458336496597, 13.2694062921357, 
    10.6859776179226, 13.9874642165191, 15.6684927432155, 10.4920141091933, 
    6.13638434279712, 7.51085197835265, 9.53300536328729, 6.754072727483, 
    3.63841916989778, 3.70434375539846, 7.71343234072064, 14.466756939713, 
    15.1680404518694, 10.8423034328218, 13.2141531523684, 18.112507400185, 
    13.7887508973064, 5.65816757080912, 5.01035326829761, 7.02398268363388, 
    3.32316079771568, 5.29614165477222, 7.43880167861388, 7.11823822249609, 
    11.5896131407498, 11.6072575645808, 10.9308422372835, 9.10646109076977,
  15.2016829712545, 15.8453332211884, 11.7969598264333, 10.5391502623447, 
    11.7424215293851, 9.9264123109634, 15.5940232709338, 15.5001785300377, 
    10.4554903596548, 17.0881509725012, 14.1908081095561, 7.30563361819615, 
    9.69213873060256, 12.5761862847442, 16.5974159481933, 15.4284350908272, 
    13.8145305042651, 14.6808266795181, 14.4171607203113, 18.45700015483, 
    18.7594727651572, 17.1719956164327, 15.0390226834691, 13.0369190416649, 
    11.0808421232646, 11.1206293158149, 15.3842754186432, 21.292033546416, 
    24.8211010739159, 24.745058239882, 18.9176823337721, 17.4855801656053, 
    20.7880547642728, 16.2179195294028, 13.3798782960964, 15.8743296090434, 
    17.3965542304212, 13.4804321349075, 6.74134792006375, 7.24669868493176, 
    13.4299708980643, 18.6408035931013, 18.439269107551, 14.3296293045992, 
    12.9774421132513, 15.3565734756243, 16.9007421631783, 13.9506243237181, 
    11.3325880707897, 12.5846171411014, 10.2289581201095, 6.02919569267434, 
    8.92599052265478, 14.0489643972405, 18.5792583871705, 16.4703751677294, 
    11.3221140086972, 9.98055055790551, 8.14703276512041, 11.3117932782513,
  14.5223903578306, 11.8335317432165, 7.79357042550972, 10.6586684129972, 
    15.7058707185659, 14.7939774593141, 13.4475511759643, 17.0143640603345, 
    14.6917502862979, 4.32727678645428, 3.54048223149461, 7.2475694487613, 
    12.2818547110066, 19.1767409896788, 16.8341591431176, 15.8125207571174, 
    15.2788498299513, 4.58725429441597, 8.9127307081281, 18.6867362894681, 
    19.0173159216242, 19.5759969722418, 18.6804796106362, 14.3965257011474, 
    6.67976744832814, 10.2926793329309, 19.1330664286291, 20.0389029400013, 
    13.4698718714749, 13.6534696665333, 18.3765529308744, 17.127035192221, 
    12.9178123149429, 12.5949023480079, 16.222626476147, 12.9479203063864, 
    14.7195266879386, 15.7051643323255, 15.2497634593964, 14.7989227176351, 
    14.4054914782037, 15.2876722462526, 17.4291012467754, 17.3979480481174, 
    15.9202015345543, 16.529814674304, 15.7697566165875, 16.2490943754899, 
    15.8928141420054, 20.5313347812997, 19.3497707322241, 14.8786004083937, 
    20.178826512754, 19.9547451198454, 16.5256343017239, 14.711375725938, 
    9.35939111412064, 7.2574075097693, 12.5117174349017, 14.678463002519,
  7.66136492038222, 1.5865040813267, 2.63707691733977, 7.82657141154766, 
    10.2293236203746, 9.65652143432505, -0.269718511970675, 
    -2.01905016989601, -3.47452852658942, -0.370073182382406, 
    9.29599180262312, 13.9805357837914, 12.5826539679265, 4.11111995127347, 
    7.8291902344165, 9.89179368142698, 0.324367819671343, 1.18503216492372, 
    16.8925555578185, 26.5173303151553, 9.95849940922003, -5.30599541943818, 
    -0.217113783401525, -1.54210862374229, 2.22558673838611, 18.343104593733, 
    18.9047900018757, 18.0165231651619, 13.0529997796499, -0.596220414964777, 
    -9.71645610586584, -4.98916329251247, 9.24203639466433, 19.1553293080842, 
    20.0509525352273, 15.3439793787547, 6.55386740805775, 2.10241981309417, 
    6.10919173223435, 10.1890559286732, 11.4355710719121, 9.43132172804127, 
    1.65973527018, -4.5058625194603, 0.963694099555292, 11.1802633347728, 
    14.3200088398142, 11.0327924651076, 10.5674084701235, 3.66384044298138, 
    0.18683970630889, 4.40525173606057, 10.1427002496082, 13.6550495437541, 
    10.4818558439526, 0.7205254724263, 0.543500070447584, 9.6561146841356, 
    14.0240773128684, 12.4105974301002,
  4.20732430557047, -0.451283112434219, -0.588106957894233, 
    -0.167031084154855, -4.0169866451674, 1.84379015431878, 2.58897826248262, 
    5.58501645354441, 11.5409147820436, 16.7011416638527, 4.34319007753336, 
    -3.32561608173537, -2.1108370226043, -6.24173636253161, 
    -9.80066554364861, -5.88888862668475, 8.85805453774208, 15.8427604856367, 
    -1.70016229279502, -6.63814984717135, 7.94680927899921, 10.3818428806302, 
    -13.0624699374583, -0.705296856430567, 13.3434679057636, 
    19.9442888882485, 7.68227144852113, 0.0247156294572804, 
    -3.46783651417368, -4.92586992101326, 0.613006775237805, 
    8.73463427561464, 8.30648025950352, -1.58075797125331, -6.31075337574711, 
    -4.33711670602812, -3.98847259022512, 0.345493338528027, 
    5.55394175751802, 12.6038314074331, 9.83914662067318, 
    -0.00968782556500429, 1.03686916847076, 5.40888853646755, 
    6.38630661704191, 2.74738087029551, -2.4687153194729, -3.65748966499854, 
    -0.153315626644052, -1.33150476079142, 2.66977247400171, 
    10.6126954527855, 11.2806337507623, 1.02742399336919, -3.93792979668757, 
    -3.41720968059237, 3.29854758988824, 5.5764776136196, 4.33679066094599, 
    7.79408788536192,
  -7.96863929795913, -1.72712268429492, 1.52709815603172, 2.90288138250867, 
    -1.7897399429149, 6.93969547337231, 8.28909491565509, 13.6247092483947, 
    -9.62135841043592, -9.82875122131726, 1.43840340344707, 1.54901064275733, 
    1.6256229473786, 3.57518871763729, 6.63958021472925, 12.8266236255107, 
    14.5608849225393, 2.83877231177107, 4.95271416782783, -1.38415621148557, 
    -8.23353545044218, 5.74576066624833, 7.78691210285684, 12.5409017163488, 
    7.13698684647456, 0.666860665364204, 3.93144965077121, 1.9284920432207, 
    -2.37159243376078, 0.770420325020968, 4.15609979604871, 2.70744723318297, 
    2.61547243303935, 4.56990586589775, 3.07279300371708, 3.7665349891566, 
    5.7174159381913, 8.5304661457659, 6.19041507502351, 2.26851569154359, 
    -0.211231966264037, 0.550844486991446, 4.20095658966853, 
    5.85028310558845, 4.64703924390743, 5.67611217829042, 6.5293519262904, 
    5.45176679487551, 4.94620731200533, 9.83417837809993, 10.0122437942057, 
    5.53704655582201, 1.28296819341875, 0.934486710805623, 2.14632436565837, 
    3.16583465450385, 4.40856115078284, 9.56260708950195, 4.55507406781763, 
    -3.93817970988411,
  -1.50868888645475, 4.41046719253643, 4.47152908749887, 6.34848777661635, 
    13.0258214921537, -1.8112927900054, 13.9880886329039, 2.66445434271092, 
    -7.81508645406657, -7.58895061849136, 2.35489788410061, 3.5560874082006, 
    3.07299094450094, 7.02834249294885, 4.59742973384281, -7.86108160650035, 
    -4.47058365327121, -3.71029976596197, 0.891239003423828, 
    -1.32021864451954, 2.06335489038803, 5.18432204568986, 4.54690486079848, 
    1.20991521469068, -1.08618400666673, 6.06670173490095, 5.68782817232506, 
    1.91633719987854, -4.28780597077813, -2.05007545701165, 
    -4.05142328026366, -3.21065967994762, 3.02280672513459, 5.7520494609958, 
    5.89893281560838, 6.67168370961823, 7.54994434755099, 2.35668238582425, 
    1.04308081857789, 1.22635680959949, -1.39970649918089, 
    -0.929807355253871, 0.107147850242043, -2.15539702665453, 
    -1.20921498232048, 4.28551780078886, 5.49646687769673, 6.81836911477802, 
    7.95972984606652, 2.39586920388362, 0.0461887049363677, 3.23206893178969, 
    -2.01675500415411, 0.499058259517903, -2.04833436060926, 
    -2.84366447342529, -0.0836759649835878, 1.85299362691444, 
    -3.86875603818617, -10.6446796873056,
  5.52542458781334, 4.41492511749755, 0.389100850124894, -5.79593104006795, 
    -8.2610251851135, -5.80856787345154, -6.02140539587025, 
    -5.81046947533686, -4.04122119068974, -2.31652382270467, 
    3.76784279479469, 2.54678611963273, 3.85928661696603, 4.79821361250489, 
    4.1730073922663, -0.262619562886405, -0.150648238507857, 
    2.39289616067029, 3.30573892652257, 0.174648672535725, 3.96737815535989, 
    0.997571206540238, 4.54690480923727, 3.77820493560327, 3.80732260858437, 
    7.7346726623828, 5.5114143471186, 4.06933955739907, -0.0586753570709367, 
    1.18556455599173, 6.65378169118994, 2.13390238456467, 2.95623168852529, 
    5.12945646243953, 5.08047128356842, 5.2831139806184, 6.06585939597289, 
    4.15409717009662, 1.03042739088992, 1.66685290958803, 5.55759510379599, 
    5.53363419996725, 8.56326208169974, 4.25354793721362, 1.60394539134953, 
    3.83735975009937, 5.98682489873596, 5.4806378486453, 3.29588274292987, 
    2.24076350203527, 3.07238624938098, 1.96191135211398, 2.09880953935839, 
    3.45006319098493, 4.623535346171, 3.3625945254102, 1.0362984820908, 
    5.10404933835313, -5.2990243491836, -5.75254720926751,
  4.8965640956652, 2.14281713934228, 5.70324237345773, 2.86931056267456, 
    5.79839446039786, 6.1999406899002, 2.89945336748994, 4.43383044328759, 
    5.3222343305223, 6.44796749082125, 6.7209260502075, 4.48306485899186, 
    4.64081902599782, 7.87323237091192, 6.37366271505225, 3.78550647681934, 
    3.30210227660549, 3.68753944061136, 4.65139220769486, 7.75416236141983, 
    5.74511049128475, 3.47256876241335, 7.61400588440113, 8.16304122910863, 
    6.65301151052644, 2.19159541582772, 0.196830811541833, 5.32381829618676, 
    8.37059265582204, 9.79918994752926, 12.1251961692852, 12.4763377608171, 
    2.33569955316039, -1.64028504073622, -3.06905956884962, 
    -2.33720333351136, -2.43711659986572, 0.962536433210695, 
    8.06919240377935, 10.2877627886439, 8.35793988432021, 10.0733707027352, 
    10.0356850879698, 4.4348834215217, 2.8014857067499, 3.12471452231018, 
    6.35837876216221, 8.54955079037972, 5.27429621950261, 2.02779228528516, 
    4.85126002104998, 6.26622892541805, 4.65609960947072, 5.62781952809296, 
    7.24830496322291, 6.11701620577706, 4.06418461943983, 5.90263361178287, 
    7.74125877870917, 2.26734435775738,
  2.23229341000941, -10.3277293634657, 4.44356780581271, 7.55045384843856, 
    0.293645469977008, -1.05997708391604, -1.37094211574635, 
    1.94775168413783, 9.05934286310463, 15.4654647925217, 12.5769230835271, 
    3.77644188876898, -0.473953758307507, 0.635023427577463, 
    5.61920430861512, 8.60417308181423, 6.47659566121136, 2.69667304123627, 
    4.87534547065873, 8.40878826902048, 7.73479408454367, 1.28637142557665, 
    1.44886721261711, 6.04390812720058, 9.02579265523048, 8.55068468543419, 
    3.83737027616476, 1.45378636293657, 4.84446310135983, 5.3223211636456, 
    3.46837206453425, 6.93833182524392, 15.7573319933326, 8.81317362328604, 
    -2.7258716790931, -6.28350656145706, -9.88234517078456, 
    -6.88159346128585, 0.916335565240485, 9.24859191351862, 10.228709934808, 
    4.23472250686292, -0.249785706246428, 0.454423642229772, 
    2.89248691488559, 3.23349732641365, 5.40652352618147, 7.93140248224988, 
    6.98855402107373, 6.67210842530103, 7.54538157651238, 0.961104704599541, 
    -3.45768587115938, -4.28228827468275, -6.28606029264864, 
    -3.01972830766691, 6.12229818669746, 15.4848962930641, 7.79574592435475, 
    11.1030516129502,
  15.8519000425583, 12.792917083902, 11.0185874199032, 15.6389322510169, 
    17.9519057044732, 12.2263546572683, 5.5518529259848, -0.186895683105778, 
    -1.42229561618205, 6.87775446319115, 15.6248213209576, 19.5257167984069, 
    13.3868337614348, 0.813457263695267, -3.53621423310771, 2.98401549550728, 
    11.2815579922054, 13.9344517280056, 11.0266032216272, 5.1823913194338, 
    1.96575117842274, 5.48193396286646, 9.74543237563295, 7.86203518375186, 
    3.2873425334652, 4.50628844934659, 13.7177540927473, 17.8365351201891, 
    14.2853627219535, 11.4322866077074, 8.34299427595825, 4.97152005488746, 
    10.8888483448528, 16.2784599210074, 14.2200497899523, 12.108344688835, 
    13.0859421383826, 13.070058110577, 9.9973785683086, 8.47715283151144, 
    10.2187451940705, 11.1507527385901, 10.384841489177, 7.94555024173623, 
    6.62712946668366, 3.76116810007997, 0.131375016673685, 4.37328811337792, 
    9.52100357669329, 7.42222187660584, 8.38340971127249, 13.1922917221245, 
    11.8575001395332, 9.36874004085075, 10.7936491175415, 8.97066933344981, 
    8.31853891160285, 13.0460827139803, 18.392378566953, 17.282697636688,
  20.0974828395137, 19.2086853101319, 14.6119484040158, 10.8919764359513, 
    9.70875572500942, 8.94824264667913, 9.91273400384737, 16.4601892590924, 
    16.829709634934, 12.9665746349184, 14.5103666058595, 17.4657666842349, 
    14.8162324760951, 9.52937959902273, 6.55528705177206, 8.26826250685178, 
    14.1641634389203, 16.1481391866945, 10.6599801967501, 5.71107944396856, 
    5.07381580277414, 2.80174245621312, 8.18132318931055, 15.9089412221733, 
    17.5762381858827, 13.4364997841538, 9.19407830423548, 10.6566226028394, 
    14.7428511395334, 13.6084696540509, 11.2647273234654, 10.9055634345866, 
    11.3260076437125, 14.7566684262138, 19.4175422753906, 22.1707086185225, 
    17.7578021163413, 10.4576243294586, 11.2707140636505, 12.9101965446912, 
    12.1648938894334, 13.9501812303652, 16.3475495227798, 16.0094977106337, 
    11.8843506538012, 12.4463321664038, 14.6383483190956, 10.7414722609165, 
    7.99408141489875, 9.58855635528245, 9.77292341704832, 11.8233510048949, 
    16.8985738356945, 18.178939431272, 17.3362992453028, 19.1600051226459, 
    21.7579088413593, 21.3083949515968, 23.0610055091712, 22.8324628238705,
  9.48828620676849, 14.4637400107266, 18.728990357331, 20.837846320873, 
    21.4830277355057, 25.6793640146597, 26.3750563638079, 16.633534240558, 
    10.2109670601582, 9.52433648086291, 9.17032678659418, 8.54112652964978, 
    10.7646125127236, 13.1867918041717, 11.9970500225353, 11.6616033250596, 
    12.0838440540184, 16.5524070402593, 19.4740377937417, 18.0784343977431, 
    14.1955576245893, 12.973274482131, 12.3105313803454, 11.2649804647139, 
    17.1217169108235, 18.5851496954338, 12.7649398739414, 8.59071782440804, 
    4.9361230398413, 6.90314642091302, 12.7315175900684, 15.6983659004759, 
    16.1674331499546, 17.3270659244746, 19.911308118056, 17.0097182870109, 
    10.5374952336441, 8.83690833020415, 9.21208678384593, 8.90636279911781, 
    9.52647786906607, 11.5281846538051, 12.6468256955482, 12.0641499738938, 
    10.0348707553396, 6.67444428910462, 6.30335147872863, 7.83038718219903, 
    9.63820623300893, 15.422830082885, 19.0791315478054, 18.686590141508, 
    15.7319640326068, 12.4340696309147, 12.578609105425, 8.80654801093557, 
    -1.52862601380648, -11.3689739727441, -13.2808444004562, -2.94380276385016,
  15.307443853068, 17.8494473551126, 15.9354643750743, 14.3052686226757, 
    14.4231729359961, 10.4246466419144, 4.39738332985754, 7.2491921503154, 
    12.719558583759, 9.52406376920879, 2.96513518521654, 1.9083009130545, 
    5.01857637876215, 8.84724511289931, 10.7083137588101, 5.83954789124472, 
    -1.85788608437231, -4.38365022431164, 1.79130812315034, 8.12489879356589, 
    10.5464599661076, 13.5095887397891, 16.2081785834811, 16.5907065944845, 
    10.554108730482, 5.4492688456129, 4.81852990827992, 1.18206928509459, 
    0.758850871270283, 2.8247309847411, 3.56546354423015, 4.88675013869724, 
    4.7467552328324, 2.70902631750886, 1.3265469711724, 1.78017508844105, 
    5.47448192489146, 10.6847710110802, 8.84880201821201, 3.85440752472226, 
    2.4200746664093, 4.90220866923599, 9.23037731418687, 8.69361460678428, 
    5.82989050784843, 4.8086814497642, 5.79021081588852, 10.4854028963106, 
    16.1231871501768, 18.4542645841819, 18.9391132091684, 18.2778680061084, 
    20.3003253606848, 22.4485802750498, 11.5323858437779, 1.35750883317158, 
    1.41834752976868, 2.8265650636633, 5.29000532176665, 9.40680540710001,
  -7.1256587850485, -10.8015073491679, -11.8647303191801, -12.8635664704553, 
    -12.9086851866561, -8.62725728428604, 1.4982754646369, 6.31463264934556, 
    1.79728562397081, -2.87545967353593, -5.36920660893667, -5.5824548171201, 
    -3.16464759317619, -1.22187379058536, 0.602220289290917, 
    4.52206844809523, 7.08128096596709, 5.40021687522642, 3.10424061334727, 
    5.81914214109324, 14.2305032485213, 16.5994890248408, 6.02961675369547, 
    -5.45881792931512, -5.66920166229356, -0.374215046270033, 
    0.686547772444443, 0.73668546907683, 1.78754646544162, 0.310583205316242, 
    -2.99998320723586, -6.83373905900011, -9.98253510727255, 
    -11.6170248146679, -10.1288668638095, -5.03380772832678, 
    0.759112899408888, 4.43954726515166, 6.0502929049959, 7.42428959942723, 
    8.63466799941919, 4.2854568370654, -3.74573686220259, -5.11362952947727, 
    -0.142256966534226, 3.71375550356324, 7.37613897475874, 10.1590258047653, 
    5.03882249994109, -2.30499038078102, -3.36334375364541, 
    -2.60951411622411, -4.26374019538653, -5.52679529097072, 
    -2.07410805174802, 2.74840567672385, 2.69622725191236, 0.743933112786799, 
    -1.01294095253099, -2.99651233887625,
  -3.50123815281885, -8.46447381237077, -10.0091385059046, -9.35538460375735, 
    -7.79495501488118, -4.13202844489336, -1.93812581772989, 
    -2.19111065523898, -3.18767918459381, -5.07427256851806, 
    -5.65813930956767, -4.49159570115592, -2.98250708009211, 
    -0.331779280562788, 3.35906662202781, 5.39741236351557, 5.62742633406877, 
    4.92924074101632, 4.32290663332552, 3.10862450013809, -1.84538291161866, 
    -7.05516632539647, -7.54654091845157, -6.61403864450592, 
    -6.01818646494174, -5.2359404831477, -2.68374545729258, 
    0.701875521339513, 1.60417162364807, 0.857494813214198, 
    -0.76728292908824, -3.92899378334658, -7.18955908735575, 
    -7.18624347191782, -3.7608736743958, -0.356838373230493, 
    3.10907978485507, 7.01684414297565, 6.65829649957991, 1.25965757744106, 
    -4.62558601776017, -8.57402964576133, -9.05675099229013, 
    -5.00247797319529, -1.17111729363608, -0.45871761919747, 
    -3.96878808199388, -13.4201756150058, -19.9567391985485, 
    -15.7115211654514, -10.635671189896, -12.1541235641345, 
    -12.0060536380323, -6.69412281596326, -0.979492633640607, 
    1.84296876820349, 2.54920168941823, 1.87752466185049, 1.55528352308872, 
    0.682973882106677,
  -0.577774339123505, 0.584139793521296, -0.100154622585892, 
    -2.17058516051182, -3.767352097622, -4.07523952952263, -3.03450333001313, 
    -1.56779896417928, -0.626132094340323, -0.461162842118259, 
    -0.3656839021424, -0.363366526919813, -0.215496923347156, 
    -0.773158763528766, -1.73611884304437, -2.10475445967657, 
    -2.13806759803974, -1.84074386778583, -2.65737714026987, 
    -5.66172193544925, -7.79183016770115, -8.42733126305469, 
    -7.98553354916196, -7.41939208946897, -6.90611158334667, 
    -5.63419836320109, -3.84043201266553, -1.99330391350459, 
    -0.12945050713802, 1.79361832876533, 3.07863418282726, 4.67594987829717, 
    7.25089127762933, 8.24586377109048, 6.19863045210929, 2.74953801710175, 
    -1.01896018330663, -2.73054501584816, -2.7042182856997, 
    -2.49971872219757, -6.47678846381662, -8.93569172471589, 
    -7.71344003084092, -6.84192277072041, -6.03331115999438, 
    -4.55133744128616, -3.08614415325683, -1.10691314139838, 
    -0.273308629710369, -3.63018008195356, -7.58364806349348, 
    -5.57267500412504, -1.66635688095802, -1.19948674960543, 
    -1.38002691412087, -0.497321621057849, 2.50454720651072, 
    4.40233139989804, 2.70348356046771, -0.891970264476327,
  1.68376751580007, 1.48524429431077, 1.19409394279438, 1.60859605020786, 
    1.83032363543927, 0.802094834065347, -1.00712608990494, -1.9832814539759, 
    -0.559819545728218, 2.0938175417096, 3.75073996179103, 3.78981970831084, 
    2.85732029323558, 1.74071218881916, 0.565014149157892, 
    -0.606194430856251, -2.22700281184719, -3.77889077373949, 
    -4.05521654228833, -3.62271745920285, -2.6709285053581, 
    -1.80434161043362, -1.55324378376374, -2.28139290852124, 
    -3.56031455203977, -4.70120322506542, -4.92891558752845, 
    -3.98069685855062, -2.2327445416836, -0.338588492292215, 
    1.61858781785341, 3.48432772140118, 4.51528026009768, 4.51436050587695, 
    4.47499619689413, 4.08862444060598, 1.51658901981008, -3.75089575764712, 
    -6.93846682808, -4.36615972444109, 0.304625106354932, 2.73542795537072, 
    3.63611130191083, 3.54981598720404, 2.24636236784234, 0.481333562749429, 
    -1.09615043210499, -1.25610660272467, 0.0745108123459688, 
    1.23297361624757, 1.38116435706659, -0.387986078947379, 
    -2.89061897946163, -3.47996281175256, -2.88473548966826, 
    -2.40705461890874, -1.53557069996854, -0.0664249784608784, 
    1.43670635727972, 1.88620857195077,
  2.17635708197351, 4.54196892456989, 6.14585209735266, 6.73575515765638, 
    6.50348780009295, 5.52173154219198, 3.92567725394207, 2.23802550847858, 
    1.26427872173754, 1.48178538720894, 2.92148668390306, 5.06365899364107, 
    7.02078705640559, 7.81159617263567, 6.88536156854899, 4.358883553022, 
    1.33169429667571, -0.60860011992179, -0.769597889291479, 
    -0.122022675434812, 0.280788424084866, 0.334350487985563, 
    0.812343471261015, 2.20349777342831, 4.19840603657901, 5.9629513452143, 
    6.70725219839719, 6.11167082013329, 4.55127485444629, 3.30756878001993, 
    2.8501358481108, 2.56056379834665, 1.6381030296012, 0.348598699708331, 
    -0.295255746146395, 0.0257818240610081, 0.417160480535477, 
    -0.0710120693400239, -0.573952018372589, -0.145142709190773, 
    2.22344948435466, 6.29776540330179, 10.2820901784304, 12.388079467429, 
    12.2342395789338, 10.5574135807546, 8.66211545870045, 7.40368251572219, 
    6.5389088726411, 5.88793565265175, 5.38284022135045, 4.30449474926694, 
    2.51631295427863, 0.837641888823681, -0.0460485664936165, 
    -0.319480992827943, -0.642635274216192, -1.20016874460557, 
    -1.16248855648483, 0.0264843796938529,
  0.74074509532215, 0.126626420191737, 0.336993964633017, 1.20305880800353, 
    2.38289106190129, 3.43968684789516, 4.02759880748413, 3.96242649449495, 
    3.20691873630555, 1.98424846246606, 0.793213850459193, 0.122539457854697, 
    0.120599234356533, 0.638857428966757, 1.45640626191787, 2.24024120911355, 
    2.99030570620097, 3.75240274442403, 4.67963414285386, 5.92703380359611, 
    7.51386836939963, 9.2226162780401, 10.8031838762745, 11.8355937381238, 
    12.0326360928029, 11.2260623155563, 9.55565296963213, 7.31788166940545, 
    4.91794538544724, 2.7714401630203, 1.18854543454831, 0.303589714473522, 
    0.210677590273362, 0.778617344574754, 1.81903110306679, 3.05403995285673, 
    4.14722378148002, 4.7220026556327, 4.91361419277323, 4.74289022797154, 
    4.27387483648438, 3.79912532653597, 3.52674942088517, 3.50052144968354, 
    3.66589004414684, 3.88630594631888, 4.15004279265587, 4.46569163069251, 
    4.81490981387037, 5.23813980898933, 5.77224709864902, 6.52422787107234, 
    7.47017350798683, 8.41306442942634, 9.04611017762794, 9.020148294755, 
    8.0332151663864, 6.20556869186457, 4.09339342555053, 2.17223923065036,
  -0.617874974941132, -0.268925558628708, 0.00788293367202502, 
    0.211703208867141, 0.348189575595237, 0.422920213401131, 
    0.432906263646322, 0.373240242027899, 0.267152404560033, 
    0.101672475390682, -0.135134077220444, -0.425263420688432, 
    -0.731064381722657, -1.02391036924992, -1.28840964000508, 
    -1.52221973585139, -1.71579900574713, -1.88088389918065, 
    -2.0194967128975, -2.14603341769393, -2.28689993797557, 
    -2.42248487564165, -2.54298006226859, -2.63623975601549, 
    -2.6889725434073, -2.65895858216735, -2.5326646165701, -2.25116385792519, 
    -1.81628461270885, -1.32172772712978, -0.886056455050266, 
    -0.559441392032026, -0.38579377172551, -0.360031528725803, 
    -0.464547392838754, -0.647103271955098, -0.868909167867164, 
    -1.07317581392372, -1.22423410542862, -1.31247039970714, 
    -1.32971565279347, -1.32000931387792, -1.33941891094273, -1.412950504012, 
    -1.54393486913907, -1.71960633359789, -1.94766078502647, 
    -2.2196008886318, -2.51449040792611, -2.83144300895434, 
    -3.10227735196771, -3.2815786853997, -3.34642500495909, 
    -3.29093116062076, -3.11070360118547, -2.78722576157284, 
    -2.41031838685094, -2.00497017484511, -1.52137805363535, -1.04150331242319,
  -10.9218631457438, -10.7369312127823, -10.275109129691, -9.49422654806073, 
    -8.39187677878739, -7.00225636967947, -5.45288836505029, 
    -3.88121827277366, -2.37372085368607, -0.961968795032772, 
    0.285078315606862, 1.29635417820733, 2.00170776893024, 2.40801318839111, 
    2.5317050410381, 2.42674054250274, 2.21940115941286, 1.94546073955659, 
    1.69120333008844, 1.53991725200172, 1.54114562358639, 1.65906308704848, 
    1.81223153522193, 1.91887627964036, 2.02345342265019, 2.11460693793019, 
    2.12051197741645, 1.98350982604807, 1.61461260260679, 1.04196674206504, 
    0.355801929476348, -0.422986119100788, -1.24598506868272, 
    -2.05792376507887, -2.81257821607567, -3.47416976220931, 
    -4.00408392680464, -4.38682320251573, -4.62216479552533, 
    -4.70805709629024, -4.63437329794206, -4.41379770458984, 
    -4.14396210000748, -3.89763058464295, -3.66719577966448, 
    -3.43881768553373, -3.2828068075815, -3.28035874300941, 
    -3.45696170602855, -3.80993539786523, -4.33914735929573, 
    -5.02540510820969, -5.83207428821588, -6.71992313262733, 
    -7.62859775809717, -8.51671516183499, -9.31638648161067, 
    -9.99043973240822, -10.5088233230456, -10.8374635435405,
  8.92095392586832, 9.81920996176802, 10.3377251748396, 10.3046647346761, 
    9.59971934179597, 8.2265516620318, 6.56597895118108, 4.98858115456455, 
    3.58161905699128, 2.15787098727599, 0.575829016331361, 
    -0.890616504543565, -1.74086639002688, -1.753897197954, 
    -1.09945226412677, -0.0495953455769627, 1.08846012124091, 
    2.20150220543985, 3.30569291579997, 3.24971303015199, 2.1354891570704, 
    1.27880608984159, 0.884964765661975, 0.739834141035783, 
    0.617604279950772, 0.386172248525655, -0.0828477105656019, 
    -0.818988961430317, -1.49804891667284, -1.82019228333358, 
    -1.73141894659009, -1.28272331245587, -0.793421811678112, 
    -0.60541751010536, -0.855395173939208, -1.43689689938044, 
    -2.08359932511225, -2.41066698884553, -2.18627313972067, 
    -1.38806326312141, -0.0944641047613717, 1.55485404963566, 
    3.32436688925477, 4.74137528894185, 5.28380593004107, 4.9313638815548, 
    4.06541345594511, 2.97528388620233, 1.94402996594397, 1.33019880515652, 
    1.32245873956147, 1.84669171843452, 2.69095889781834, 3.59032317317167, 
    4.40679030300417, 5.09106553133165, 5.56150095976975, 5.98311640117681, 
    6.72161957681992, 7.79630137556583,
  3.5188719742317, 1.9405541067585, -0.338352495956148, -2.11304366672807, 
    -2.2879469995264, -1.32227592787478, -1.16486207508914, 
    -3.11519873016916, -6.12504452031783, -7.7849857078128, 
    -6.58591594565726, -3.15518430638054, 0.204095275999539, 
    2.49585256728803, 3.76890860105334, 4.2731063467322, 2.64233835451215, 
    -2.01121943545715, -6.98319076519645, -9.89676309407795, 
    -10.0616434376053, -8.36789135584157, -7.01742712274998, 
    -6.04973981868205, -4.8601066418879, -3.3964134460013, -1.99718526350309, 
    -1.29529653937341, -0.858672918798681, 0.42260138252629, 
    2.77450593937625, 5.18056177896437, 5.92801946326097, 5.03972026352123, 
    4.00181217701051, 3.81577936736592, 4.62561026033665, 5.7700987817594, 
    5.70279667039741, 4.40166572687507, 3.39503660877563, 3.04287486771526, 
    2.93206366096524, 2.9832851009622, 2.73512575801793, 1.94131788574325, 
    1.30536759828862, 1.62392243405677, 2.99583471163324, 4.39041024450504, 
    4.49405974433507, 3.59189510012583, 2.72406466092213, 2.3111893856287, 
    2.35468798333576, 2.85457095819496, 3.30954083031711, 3.99437664702326, 
    4.43927152502966, 4.26053808022147,
  0.960170709241924, -0.581455952431253, -1.14156453217558, 
    0.335856849188174, 1.35056656448155, -0.952428392138106, -4.852499303133, 
    -7.31729449018119, -7.5937377927289, -6.8988941368351, -5.33793087970133, 
    -2.88667361116438, -0.22298105188955, 1.44982823215551, 
    -0.0352413890295661, -4.14660124931058, -8.00765539674943, 
    -8.33964494560825, -4.05846926636141, 1.29303616445135, 4.0472012369803, 
    5.64616024443543, 5.66647009328254, 4.24901008652514, 2.34355517865423, 
    0.370102634454206, -1.30656466279734, -0.330742851248915, 
    4.73405416167477, 7.74669319652271, 3.37049298895344, -2.09161100179761, 
    -2.28836761336452, 0.63754839401961, 3.32705502161852, 4.97494681187082, 
    4.57639227235386, 1.78436923825059, -0.20876394382912, 0.921727460816063, 
    3.30671321833897, 4.199866531414, 3.33751274641995, 1.76581686458858, 
    -0.208783264603452, -1.47585048956137, -1.00395471765106, 
    -1.27138023795358, -4.80061801659498, -9.0652834884104, 
    -9.79223667644394, -5.83687455288705, -0.397438197492432, 
    2.32995182965486, 3.32185701365162, 4.22838554120196, 2.48954334836509, 
    -0.632427721064592, -0.939456627044507, 0.711628740127867,
  0.319753038271723, 2.59095510043389, 4.01800943566186, 2.74813275959893, 
    -0.848219327491182, -2.00180554874973, -1.19369298866755, 
    -2.93052168412851, -6.96713077544143, -9.47017942810067, 
    -10.8301879272906, -12.014635000089, -10.2700499782953, 
    -7.99794119802943, -7.66149620808957, -7.50867583581704, 
    -5.72577551461056, -2.4371478473391, 0.332148897905576, 
    -0.908703811259549, -0.0391668766979617, 4.40455459759163, 
    7.78270811632487, 6.15626626761613, 3.33432352556069, 1.29451620929508, 
    3.28198642480026, 5.54147355520734, -1.10105795645554, -9.44617549289352, 
    -7.31177063163252, -1.24997400522963, 0.384542869907902, 
    0.483536009838085, 1.14760240358785, -0.500998340687753, 
    -2.88464391027215, -1.82115636035012, 2.32603470330195, 3.4845396230723, 
    1.41595436304661, -0.740943573011996, -3.12006206096312, 
    -5.03045136936689, -5.17010667184319, -4.20527158040812, 
    -3.6271543861824, -3.20070237350491, -1.67413535450771, 1.14511612767738, 
    4.17977255961583, 5.65288919393178, 4.86186832978252, 4.05861501335509, 
    2.04103812284188, -2.64077686652066, -3.45517806449436, 
    0.680775952420139, 3.07395481333396, 1.24877591213366,
  -9.40914784730576, -7.18317113447224, -7.09812692590924, -8.29964019963946, 
    -7.53115367494229, -5.61002335702066, -2.49379330146684, 
    2.35950907214378, 3.47670518260636, -1.15911219988912, -5.81545948700167, 
    -8.52574171709291, -11.5029598801138, -8.22303788072418, 
    -5.05586722525417, -5.06771200306788, -3.06008713070168, 
    -3.22161935522872, -8.33258604060759, -11.2807258006506, 
    -10.4483529546934, -9.16532018169839, -5.70582562601846, 
    -0.768277537208746, 2.95530970801572, 5.24845306283818, 4.38513508978322, 
    -2.92149343267345, -8.07254754430104, -6.04684181340395, 
    -4.20490474394804, -2.53274488427538, 0.608076489633496, 
    0.312979512784771, -3.20856263760587, -5.6182526527156, -5.1320488070812, 
    -5.56222737721811, -8.03911559536713, -8.11976688050517, 
    -6.87714789073019, -6.65377106870291, -6.26166340643877, 
    -5.85614083851571, -5.55588206294827, -5.37985046789404, 
    -5.36893621527482, -3.98327986763029, -0.24554613300674, 
    1.11660271478145, -4.72112469059169, -11.1876427578187, 
    -8.76249024212859, -5.26828877424649, -6.71220080108077, 
    -9.01647113157375, -12.0330594070973, -15.8449818590909, 
    -15.7121343578743, -12.1738895930583,
  -17.0740158068013, -14.2361588217459, -6.63974220019966, -1.97846262366239, 
    -0.482498829835768, -0.105800377721861, 0.125469322973244, 
    2.28400275122046, 7.85213517591353, 11.8108893080158, 9.68316549088029, 
    7.80294257243689, 1.36445582877127, -11.5346266756298, -7.42550452246976, 
    3.08052658049809, 2.73501473529241, -2.40567363217125, -10.2791858699122, 
    -14.9160603689776, -17.2670192498275, -17.3644026546194, 
    -12.4340717283167, -7.48792647516575, -4.9028404520681, 
    -3.24126086169154, -4.22999078521192, -5.20961936698179, 
    -4.20760396915826, -5.4960407232196, -9.54554905934003, 
    -13.6130293608726, -14.7555458917701, -12.4585940095952, 
    -9.71715835296572, -4.69128026702124, -0.034818760903288, 
    0.900009703575718, -2.23520196972134, -9.18493158291756, 
    -13.3831343757364, -11.8744136813426, -9.07137482011506, 
    -7.75240715985451, -8.70446843124393, -11.0144539145377, 
    -12.9313852180154, -12.3678339704521, -7.67983610505107, 
    -1.05353928958389, 3.64333302546996, -0.419261237007176, 
    -11.9172836617843, -10.8847691588724, -1.43410464494397, 
    3.63560813514937, 6.70409144342622, 7.39903108681156, 1.54542981374907, 
    -10.1251043965052,
  10.5173949647137, 8.39201058624198, 4.24940024310774, 1.36504755193479, 
    -2.27548666359553, -4.79611206432109, -4.89075483028635, 
    -0.205705418983136, 7.00151771239899, 12.3363108866712, 13.125662250666, 
    7.83476769554997, 9.57650331313401, 7.48312377785578, -7.67223765950733, 
    -7.23464306532167, 3.80880783349867, 9.32478137384568, 14.1693183699125, 
    12.6514411107421, 4.10189325845903, -5.98932538349667, -13.3098758905903, 
    -11.89076084121, -10.1252264431843, -12.9227766891764, -14.5983118542993, 
    -11.2659217777332, -3.51108561781535, 4.85450435962955, 5.69886532705473, 
    -4.73758296061796, -17.2415094449367, -20.737823612943, 
    -16.4392162795278, -11.8523032845964, -5.08379614445795, 
    0.863027613035757, 4.24839909976734, 5.64259447234381, 1.5123791815502, 
    -4.67121941066283, -6.34483167376727, -4.65318095072913, 
    -2.01508468032009, -0.353210235638488, -0.925708930250974, 
    -3.99835782812029, -7.77103348839612, -4.27343037498788, 
    2.19063744043456, 5.45155481442249, 0.499870051921301, -16.9578045223012, 
    -17.8499458110038, -1.58565114840361, 6.18772831767156, 6.93040515123047, 
    4.87495582408588, 6.37183793777209,
  -3.22953372227753, -0.515647706875399, 3.60672443716552, 2.47598408732549, 
    4.61593131040952, 8.13654041791669, 6.40611803993621, 3.36310299710275, 
    1.41265215736929, 0.0222784722389546, 6.08943875244162, 12.8156898903245, 
    9.93475957692745, 7.60278767680616, 7.55677859880558, -0.520278823187869, 
    1.07229870431475, 10.9556676696618, 11.7410803228951, 12.0298111455057, 
    18.8747561681316, 21.4078826616769, 11.1196438893103, -1.90539721806627, 
    -5.63212093209767, -5.45377442027293, -8.8478316070081, 
    -9.64980093743067, -6.95936154865365, -3.74692881041501, 6.9596750171973, 
    13.7052307473597, 12.2674458429392, 16.6096126824938, 18.1449161060908, 
    8.17379364882519, -2.14691235061525, -1.61875460040625, 2.7696908457442, 
    1.6695334871919, -1.5067296790245, -3.03606073722207, 0.799697577995564, 
    10.6242351259579, 14.5902091330337, 8.94533918892616, 10.9685287019342, 
    20.233105322477, 14.9287881825323, 0.973226781343964, -1.8331894820266, 
    1.52021202168367, 0.224908422738168, 3.47285352329294, 0.992395795074122, 
    -4.45859483689629, 1.75043984969237, 4.51696428211964, 5.164561756437, 
    2.54202087223494,
  10.0077669812836, 5.79534634890863, -0.64650068406385, 3.06540798189663, 
    3.88080686713918, -0.409031328833702, 7.83757522510259, 6.82356066984551, 
    -0.0396843923605434, 11.0130346553028, 9.85604688350682, 
    -2.0909142166613, -3.77152986364406, 0.516415204078736, 9.75122337947217, 
    9.31567774886932, 4.2033051218564, 4.79071320327416, 11.7100736562074, 
    13.4404346573735, 3.67838681253022, -2.51576579539572, 2.34321585533193, 
    6.3324398962579, 5.2000329531644, 8.60412934589498, 15.1597629481551, 
    19.729486148755, 22.5888558472149, 17.0329786677184, 3.58681076374854, 
    4.80207658586641, 15.1128331127765, 9.93753658588619, -0.474774815276985, 
    6.40642241492361, 11.1340570703831, 3.92414905307871, -1.0626496507048, 
    3.07371594470398, 9.91279366500106, 13.6689004682668, 10.5202233180128, 
    2.61255706472738, 2.16530510539896, 12.2993125260831, 14.1612076702461, 
    3.67963823753785, 3.27315190947508, 4.67965815087361, 
    -0.0901271976391772, -0.401337950365015, 8.16783884703024, 
    13.8658212540085, 14.2131730763022, 7.20483089249758, -1.08905266796181, 
    0.0770339015037881, 1.73542586109529, 5.6365011188858,
  8.68630068237001, -1.96206980655814, -7.02391863442779, 1.68692618368296, 
    8.586558036926, 9.56969784888694, 6.25184341324211, 11.6707343058038, 
    15.2895972675998, -0.119328345367124, -7.39090676707975, 
    -4.5991457386941, -2.12794442320789, 7.33835414727787, 11.108366660571, 
    11.3554090932242, 4.9125757127885, -2.91773047780467, -6.44810281741814, 
    -4.10047092943447, 8.75073113092331, 15.3423053344474, 14.5259349729848, 
    8.66752955724242, 3.50562085172099, 7.09857503720631, 8.16606175272335, 
    2.48478296338317, 1.75257813685657, 6.22295834554452, 7.82364972933393, 
    9.59729905374958, 7.58368863731322, 2.44690973216584, 1.26889367049666, 
    3.79478590350133, 5.86679433059255, 1.90440243581138, 2.87804743548668, 
    5.28446683497388, 6.26610694551579, 9.62332169148297, 7.90048905427904, 
    3.61402558407964, 6.37829077420632, 8.16147215368408, 0.934597104651494, 
    -1.39077522844215, 8.166285833546, 12.1434237955917, 6.25857184584522, 
    6.77307585663987, 10.7480767983599, 11.113028789291, 5.3946940586683, 
    -1.88501147762624, -5.43348116003733, -2.68878330471, 4.25134331730217, 
    7.64628968096497,
  -2.48191024744104, -7.37523805033581, -5.09613724004093, 2.32819494727592, 
    5.21050848070042, 4.74387137707719, -0.750288056685196, 
    -11.5246322453555, -13.0201521796987, -5.43682216649967, 
    0.46770600349819, 3.74917761585823, 5.41590215956631, 2.05227909111934, 
    3.01710850399608, -2.63366717392164, -11.4417593387084, 
    -7.35542052234965, 0.317853509468044, 6.69566624097626, 3.67355763901876, 
    -5.61214406882288, -7.67543974054811, -9.44604918459577, 
    -3.39413420852426, 0.812029449597397, 8.66623398939792, 16.530565308613, 
    4.98375972009319, -9.75472527616942, -12.9557183587651, -8.9117978223224, 
    -1.07917698408412, 7.45250332465206, 12.0578839066926, 9.69300494953011, 
    -1.32996540495131, -5.22444070086108, -0.556035191761357, 
    3.36375883670057, 4.92315591033064, -0.303659545426741, 
    -7.51813348358116, -10.1347424987927, -5.52801840766677, 
    0.324231589764378, 3.50884500558014, 4.61653206991574, 2.88420027143253, 
    -7.02212618192537, -8.03384592019891, -2.23240530030304, 
    1.69135163077654, 7.40324871327372, 5.59011280632781, -5.05961986793856, 
    -7.28966614595471, -1.11837708086399, 4.0856714578504, 2.02670924448215,
  2.05807327680882, -4.78328369478953, -3.72452796083539, -3.01262058398481, 
    -6.1742190052773, -3.76569392549273, -0.521823398526906, 
    -3.40131578144719, -2.55429371073025, 3.7867740093839, 0.454754249177526, 
    -4.62764672610026, -7.76355570129971, -8.7587309219242, -11.141675196624, 
    -9.32761189295595, -5.64037661138884, -2.13992650527689, 
    -4.2138474760867, -2.71812913678298, -1.69407556077374, 
    -7.98888493410059, -18.0750545281328, -10.0826462554855, 
    -1.46994431604947, 3.83610130053029, 0.526317619778401, 
    -4.79989889121615, -6.74811387673662, -8.42144728124183, 
    -7.67974147383634, -3.2210634869508, 1.14010048986962, -2.25781260010802, 
    -5.48434038817855, -4.5145667366043, -7.17695039675587, 
    -6.59407244867635, -2.76708040643655, 2.56164827660148, 1.58792524613986, 
    -5.19830679313111, -6.89959876479857, -5.47995127933723, 
    -3.72594041622924, -2.10564865709688, -4.4650224444276, 
    -3.22698253229826, -2.60838436157351, -5.99463853224962, 
    -4.74320596292257, 0.92558765315882, 6.06752108910355, 
    -0.359184807606225, -8.64378568310319, -8.31182677621017, 
    -7.13099935277208, -3.19113236986014, 2.28476369765199, 6.64724588521408,
  -3.08509585457126, -3.88791102974484, -4.8972291794823, -4.46359695669442, 
    -3.67002531025328, -6.53912520380076, -5.38595915132408, 
    -7.02044428999033, -2.79677532785943, -4.77249402375071, 
    -3.72526247062777, -4.74705641027387, -5.04904335988433, 
    -6.52741707357651, -8.57118955461167, -11.4982440236793, 
    -9.06094393872152, -3.413273458209, -0.720016461062599, 
    -7.10568452273524, -8.10989624129715, -2.68436073552833, 
    -7.75070047323567, -6.89169100167523, -2.77373913571697, 
    -0.598260783439671, -0.501857627476401, -4.28899271853858, 
    -3.87236722012509, -2.56076349095093, -3.08402833875359, 
    -3.18788575429758, -1.68023319664624, -0.170238084175848, 
    -1.14939148207675, -2.02801506548571, -4.75375608241402, 
    -5.57205420122429, -2.40586192873467, 0.324077147615068, 
    -1.58640824294161, -4.53852070418921, -6.51155691715573, 
    -5.23478181659702, -3.88515835505749, -2.86533641525143, 
    -1.62949485915494, -2.16231258002235, -3.61299524180348, 
    -5.12975333230179, -3.42330202726508, 2.22861296576149, 
    -0.284534426348658, -0.00148881053745584, -2.64390210851687, 
    -4.45395056970446, -3.89635282985305, -1.95681651734484, 
    0.828197456977311, -2.86418104582288,
  0.0892054859767563, -6.38336595572229, -6.3426275904529, -1.45904346091811, 
    -3.55937540048609, -1.35913673799619, -5.84966932846276, 
    -2.28292673256525, 7.36908417515403, 14.4920450425133, 
    -0.627377176010984, -4.2245399505684, -3.91420624413591, 
    -3.42434066386317, -4.30073496183581, 0.108744886562905, 
    -0.71110273487885, 3.7388796005592, -1.39548119644932, 3.23728538135941, 
    -1.63334725595615, 1.68870079928038, 1.32742233934425, 1.10605554296482, 
    1.50920586346248, -1.30542959869829, -1.00137672204276, 
    -2.74198813803648, -0.873820848093319, 0.27937211224654, 3.6560780784487, 
    10.9797471084134, 9.91782357226344, 3.6840217453903, -0.772405732019556, 
    -0.992616198735269, -1.17228059594062, 0.584227894075812, 
    1.12989424020099, 1.68996637502275, 1.57754151083115, 2.43926058887989, 
    -1.22006264281246, 2.16003678281005, 5.50637203991038, 1.20460375636631, 
    0.825524620728326, 1.20977717034658, -0.4397718158213, -1.65071936360868, 
    3.89212855108214, 1.04610472258539, 4.52827693100543, 
    -0.0328938373634474, -1.0706951893977, -0.946840395741947, 
    -2.26670025904464, -5.21527563330259, -0.348108249740484, 1.14032696121377,
  2.27978109747451, 0.722882044057166, -0.764988344403533, 
    -0.391634874341034, -1.02764503111887, -2.51438792974342, 
    -5.80413005025785, 5.71598167118113, 9.12444490255603, 7.90701228392561, 
    0.969407695779431, -0.928000306965919, 1.40664495247136, 
    2.72171122489311, 2.75610185297428, 3.75125565471207, 1.19409554330224, 
    -1.64381369385372, -1.38156579457782, -2.30302804442802, 
    0.560967220909941, 0.552196312530393, -0.391916220904225, 
    -0.0864803179175451, -5.08174042449281, -3.1040893433849, 
    -4.35918674338413, -6.92378203367722, -7.61360079733845, 
    -6.89095128121671, -1.91412545399881, 0.321079141594359, 
    1.66377224693753, -1.04358235865492, -0.766995549055602, 
    -1.24579286604199, -2.67732644684527, -3.08312504873656, 
    -2.97413219094475, -1.86251056173125, 1.11905384824044, 
    0.206748383821478, -2.380549118704, -2.57929845477194, -3.06406488489308, 
    -1.05869025975996, 0.15466450064127, 2.43050153306106, 1.7636076737304, 
    1.46518276690056, -2.83570508412045, -2.13806138670989, 
    -1.49202131603414, -1.35271754916952, -1.64100588677422, 
    -1.51378625198105, -1.36494358409898, -3.09814897094765, 
    -7.97668325335114, -11.4094411656573,
  -1.04836531313057, -3.47769654248346, -3.21354521169283, 0.22410426006601, 
    1.53493803591292, -2.15585751809226, -4.6032211534307, -8.24402776781422, 
    -6.01698420545627, 1.09873824473676, 3.51415722419243, -1.99560929656962, 
    -2.35565603608372, 1.14886616704928, 2.15245036495678, 
    -0.456881688413078, -2.31848890207787, -1.73916979860713, 
    -0.372524149822538, 0.311154478493821, -2.29007464458168, 
    -3.24281307065587, 0.717162598276328, 1.30218966587369, 
    -0.0320447331843782, -3.11252909222402, -4.67952411711062, 
    -3.84818423100477, -4.73907570373799, -5.36546272911295, 
    -4.48422757503198, -1.48605564342844, -2.93048960557812, 
    -5.63620103079531, -5.12634255218508, -8.80504641442633, 
    -9.93958617896078, -8.62651699985545, -4.62331263005655, 
    -0.271663009378169, 1.69614612996389, 2.19180356019154, 
    0.596270353892643, -3.3847545419227, -5.42580105613929, 
    -4.39206414189845, -1.16112062228147, 0.592473535730694, 
    0.118615932140025, -2.13248870782111, -1.655676519724, -1.28287348716621, 
    -1.9356797543454, -3.6669699271657, -5.18768620166327, -6.16233169365523, 
    -4.27910107599162, 3.53433292611879, 1.56687968540295, -3.89006651128303,
  -11.9838615773806, -14.734581229464, -3.89528147638378, 2.44143809982234, 
    -2.47374930104312, -5.60347304196167, -9.55886233579703, 
    -9.95790714835071, -6.40515884975126, -0.138539000611652, 
    3.94050236300362, -2.82581085405055, -5.57371394487981, 
    -3.99135797159862, -3.47317533675191, -3.18610526541296, 
    -2.06407593919392, -2.6889617227715, -0.412576516834165, 
    0.232282975614043, -3.7487323471034, -8.44978874585842, 
    -4.56966625254101, -0.655103562059561, -0.572077970856068, 
    -0.68653230845969, -2.40092890865855, -3.66909167287412, 
    -4.99489966918094, -7.61828660273999, -9.93403254170096, 
    -6.6066480736007, 0.17665227333383, 2.70423153914465, -0.659341900080174, 
    -6.75724342631893, -8.87004863488641, -9.19390481179836, 
    -6.73331273418739, -0.860404539056764, 2.16503757192169, 
    -0.863239577345201, -4.04226116823091, -4.9386428626327, 
    -5.14066759707265, -6.52074295284827, -5.80937227604864, 
    -2.40227820411725, -3.52177341133984, -4.73155445520697, 
    -2.94196652055708, -4.46549721861435, -6.44911905595304, 
    -8.09213947544877, -10.4426253466113, -11.1836568711588, 
    -6.68501324887358, 1.66905489800827, 1.74893660517976, -4.27130809513379,
  6.01918903304431, -5.92083639252521, -6.46988353248588, 2.89445420488996, 
    11.9287004649166, 5.40922317418191, -4.40929298808239, -8.92056991091795, 
    -7.57493215179287, -2.34563445322575, 6.03382597805042, 11.8504169205471, 
    5.91268099596847, -7.03404620151334, -13.030516389917, -8.63962526440211, 
    -0.464089900213357, 5.53420302813548, 4.80313365383896, 
    -1.21904575271169, -8.67194281594986, -9.40035479887671, 
    -4.37666672455407, -0.172217076919119, -3.50090885313266, 
    -2.22570310161449, 7.60953320869225, 13.5399298339142, 11.7472784434345, 
    5.88350932231475, 0.461609107157381, -3.02942422590434, 
    -2.06249730974139, 3.21197050812708, 5.50052632385471, 8.87764120996721, 
    12.2141219300671, 11.0043137594404, 4.98786844551038, -0.538431701155129, 
    -1.70164136939701, 0.437894057833241, 3.53342573969832, 3.07167186731259, 
    2.40573530858057, -0.979872044697621, -6.78995886612381, 
    -6.35219471495637, -5.43486331153069, -11.2948827267188, 
    -8.94206751451604, 0.758573152916447, 5.57910340638137, 6.95699811145284, 
    7.62431564081984, 4.86897815689228, 3.39833026501486, 5.44132508902764, 
    9.39527272867926, 12.5321286449896,
  2.46953302574272, 6.26471070887274, 7.77145720244387, 1.01100611360597, 
    -2.67152121778797, -1.34165729492241, 4.30213799325813, 11.5400669276005, 
    11.6625831344869, 9.72644523770143, 8.5539555511318, 10.6400352684891, 
    7.00021547295664, -2.38064098166124, -4.96133888476667, 
    0.107708601918972, 5.96856838854066, 3.40137456982585, -1.14986738302943, 
    -3.57636277535358, -6.94009485070567, -10.234503324726, 
    -4.54190069194063, 5.76744986791175, 7.313281277943, 2.5457383183782, 
    1.36806506335469, 6.76718288449329, 12.0457948397442, 9.98657199231423, 
    8.14419493847369, 8.30091272317594, 7.13605922152933, 4.82056083957967, 
    6.44836286621531, 11.4098111000592, 4.73613611983044, -4.61056408260763, 
    1.24747632520968, 8.6860816222929, 6.75126703185185, 3.17715737943952, 
    5.83352020247993, 7.08656817541049, 3.08831602637356, 6.44771430951278, 
    11.0767845990287, 6.72616236287605, 2.36315646814266, -2.41620783603695, 
    -7.71936100533511, -4.57905243442814, 4.49952666389575, 6.45601703136998, 
    8.52816943034751, 11.1827348416814, 12.3522380365785, 20.6595069238273, 
    25.3332925675115, 15.0260589610203,
  1.6970985512445, 9.84057113716788, 15.813799472287, 18.1823224164967, 
    14.8520187642671, 19.390204725791, 20.8913147294868, 8.8144306867889, 
    4.24442455459281, 9.67771386964257, 11.3970423192585, 6.62598297367308, 
    6.90250182336577, 10.5911227788449, 6.19611944414035, 3.57225255527583, 
    9.83136206869165, 18.770995673157, 20.5355186476376, 14.6605545961437, 
    8.74169807989293, 5.09433609700413, 3.80435228191952, 3.56756219921257, 
    9.17054700794487, 11.9042710025631, 8.13377352051063, 2.27855114431166, 
    -5.03595792836355, -1.49874290645611, 7.19076499537085, 11.4153373774446, 
    15.0198755772064, 19.0290977235842, 18.6483027562348, 11.5848672346928, 
    2.42444797821603, -0.421672619119104, 2.1385108236807, 4.23820897341091, 
    5.4198775990655, 8.07005698016458, 7.70881068921608, 6.16589964863731, 
    3.99044571927592, -2.06311231521189, -4.45907935138094, 
    -2.75090710570595, 2.81280129872465, 10.489659813349, 16.3263713015969, 
    16.1552159870968, 5.61370029975193, -5.28401476647001, 
    -0.112206582649834, -2.47316730958202, -14.6989959447101, 
    -22.6598503614804, -23.8004646417735, -12.6489047631169,
  13.0441463649755, 20.4585880193643, 19.6442438355869, 18.9392649173157, 
    18.4362095884032, 8.44598604130932, -3.92331421200223, 
    -0.757818637578272, 8.559927358017, 9.09647922713535, 4.96753030655754, 
    1.33603659098795, -0.489303248016238, 1.7108641448774, 1.92228338423616, 
    -3.38794719418952, -9.20965933672542, -11.6732668411619, 
    -6.52547625839437, 2.24122710618017, 7.43497067312782, 11.6219244333182, 
    19.542386090545, 22.258427054425, 12.8357727049474, 4.65375521852819, 
    1.53714007166192, -5.24217414058039, -5.03529937310641, 
    -1.56310806271074, -0.149459251849831, 4.34087812039357, 
    6.59081619570573, 2.66878485775745, -3.40091953087506, -7.35903149288385, 
    -5.77836524005706, -0.356470143937239, 0.231909027439761, 
    -1.34567343119705, 1.22196354219123, 6.04028589561867, 11.0204195044207, 
    7.77713210211811, -2.28633685280875, -4.69402687517937, 
    -0.721694195529498, 6.42052550968546, 14.6023752652764, 17.5445959850257, 
    18.580099668106, 17.20959973139, 19.3227665996453, 22.1044005813734, 
    9.31271265206671, -2.28648638655898, -1.14418356200385, 
    -0.173414495671235, -0.538796600333396, 2.70414378492967,
  -6.06578293100348, -13.9899179313569, -17.6067503486467, -18.9887632935728, 
    -19.3488655398871, -15.9205435781149, -5.07551297029189, 
    3.09487119920148, 1.25638086380034, -4.8034392201435, -10.8558355906323, 
    -13.8213068957376, -12.5257774949782, -9.57509190072909, 
    -5.5405610006837, 1.21140162782642, 3.85325111616149, -0.273575940108242, 
    -3.39401856779426, -1.00893917832994, 7.24462667879837, 14.3589131851075, 
    8.54832566768371, -4.16556970972851, -6.25908594036623, 
    -3.07891384586336, -4.84212177997368, -5.81393532872334, 
    -4.58299766999092, -5.66497123858745, -8.51838748208356, 
    -13.2851990827308, -17.9317462242254, -20.3752584312805, 
    -20.460249524598, -16.9656909262779, -10.115395968471, -2.44030076352799, 
    3.86564488897072, 7.51108424069715, 10.5887818009978, 5.81835604605528, 
    -7.03375653970108, -12.6548568865121, -7.91507498839778, 
    -1.22382711207974, 6.41561100952169, 14.3314197153879, 11.3921814377273, 
    3.15878972070798, 0.398722177659595, 0.695690116247102, 
    -1.63852736757449, -4.79598583620713, -4.43284029250397, 
    -0.813389583723338, -1.12593283777612, -2.42221334457319, 
    -1.23021595564846, -0.552092811220131,
  -4.74874796052515, -10.8588368098933, -13.4244462757404, -13.7271670819357, 
    -12.5307574087562, -8.63298696196918, -5.18227742077883, 
    -3.76709478790114, -4.63034407963895, -7.44095300011381, 
    -9.09114296852891, -8.60280867978359, -7.15235482083272, 
    -4.10309540036315, 0.176228706452208, 3.28592971264337, 4.83825261348971, 
    5.4106511487437, 4.89720381977815, 4.63778242073434, 1.35224933471031, 
    -4.93813201318957, -9.24426367699551, -11.1861984433661, 
    -11.1625118941119, -10.627153484065, -7.67336310200415, 
    -2.69757530805488, -0.106161117952248, -0.0492709585783729, 
    -1.46206675774597, -4.65190920265198, -7.87838003391024, 
    -9.11020339077504, -7.04250697395591, -3.82194763801494, 
    0.557805700234843, 5.54690487345831, 6.41359522247166, 1.83565780767122, 
    -5.74274916897737, -12.6591349175288, -15.3771362121531, 
    -10.4079859388041, -4.05184410927389, -0.44202918208833, 
    -1.51095200174036, -12.8337814434671, -23.6237758981634, 
    -19.573234487039, -14.6594400598635, -16.5514983874452, 
    -15.9688150863212, -10.6494425283222, -5.05461945861969, 
    -1.49815160468308, -0.338021806059386, -0.726971210926179, 
    -0.505491434520156, -0.68476071275639,
  -1.94512254738486, -1.09035337891472, -2.46481615453224, -5.06029700242987, 
    -7.14720413776485, -8.12127046107064, -7.31420437458386, 
    -5.37726558564825, -3.43032121803096, -2.283415401699, -2.01555309332686, 
    -2.11529864900979, -1.9195324632307, -2.27082060401765, 
    -1.91398913884303, -1.12903021979566, -1.15513329432082, 
    -1.22666094157721, -2.70834313295968, -6.72705169727575, 
    -10.6334179627813, -11.9405982474293, -12.2964622450662, 
    -11.6013708091112, -10.8275340679061, -9.00835003428388, 
    -6.34023279478828, -4.17480112342328, -2.44111192310684, 
    -0.748042040138582, 0.636292083238021, 2.38970415872181, 
    4.75889960591398, 7.25138736968354, 6.6853286019054, 3.0870250958825, 
    0.933607937800742, 0.140966017259589, 0.218410339924256, 
    -0.867506089407309, -6.8099139311528, -10.7110360459788, 
    -8.49766704732364, -5.97221714540101, -4.37723998691748, 
    -5.01291995397775, -6.24849292632768, -4.30530589232024, 
    -2.83593020803991, -7.20538091239209, -10.821207272511, 
    -9.11990951771947, -6.21499873195414, -4.87042438570547, 
    -4.49105723491383, -3.03401834326019, -0.926222553995652, 1.34792205568, 
    0.648018604040194, -1.75416869270298,
  -2.3351519132539, -2.24852093901926, -1.19561951032911, 0.3236470870564, 
    0.654523962737256, -1.28085323376569, -4.35420022918187, 
    -6.63277063335083, -6.22712423875902, -3.01690548194392, 
    0.408309270114059, 1.64206366996319, 1.396656169277, 1.28412249919374, 
    0.71534979404252, -0.809750193497776, -2.38208482162419, 
    -3.28664734954217, -3.75759305253767, -4.0218180253248, 
    -3.79478590450467, -2.99820811009025, -2.32675475668179, 
    -2.34085658657512, -2.63095855203182, -2.75713126698817, 
    -2.40750156466187, -1.99306145167925, -1.6283473814633, 
    -1.27205137181152, -0.741554151672724, -0.065986380131608, 
    0.945404920037887, 2.18641468323346, 3.01545478596073, 2.14285178956683, 
    -2.20153883027787, -8.36818562751149, -10.8822215860659, -7.499759794559, 
    -1.46162382226234, 1.64733499304586, 2.66684916779378, 2.7765671801766, 
    2.56827256763826, 2.74126735340441, 0.83100039645924, -3.29761585453908, 
    -5.43427835213848, -3.69667106621815, -2.24246306715202, 
    -3.32977624296256, -5.74280945871061, -7.34923560245291, 
    -7.81561032197374, -7.85606943349135, -7.02186597512363, 
    -5.14592652381486, -3.27364829378418, -2.29573227043187,
  -0.735103663504091, 0.731447427731985, 2.29723615409592, 3.3095660323407, 
    3.80881030422209, 3.97402297295414, 3.51495648874811, 1.90521714539927, 
    -0.496467568245589, -2.13385399245964, -1.60903469326196, 
    0.785394306429089, 3.29012414091341, 4.15079195220252, 2.90962422825421, 
    0.493695986791239, -2.01053840678873, -3.80109552427929, 
    -4.09797892775365, -3.13035809210998, -1.77996834572599, 
    -0.698703523128442, 0.128039908682032, 1.29864653471352, 
    2.97613209595448, 4.74664638125951, 5.81594324441778, 6.01130225227613, 
    5.43519089410258, 4.65567430675534, 4.02816090142231, 3.14367164175002, 
    1.37540576220146, -0.908618082784871, -2.20888569596106, 
    -1.22221525727046, 0.682871899555499, 0.791764315000118, 
    -2.70944671944504, -6.50226242390418, -5.51221514879629, 
    -0.696750634924187, 4.03513357656038, 6.10300673284083, 5.89338433959184, 
    5.01641798187222, 4.6315850243732, 5.23783390094008, 6.34892809895195, 
    6.32134777840914, 5.45691477126913, 4.7658257561804, 4.28554148411927, 
    3.53684846661978, 2.60436055785291, 1.76475059690171, 0.913826921404431, 
    -0.20253353514725, -1.27936520621476, -1.55918794531986,
  0.560074746318455, -1.18272815236122, -2.27979166650581, -2.38463247908161, 
    -1.37043405001188, 0.511276190920316, 2.58007572571746, 4.08332254245442, 
    4.53761166054559, 3.87612996743651, 2.3412133586789, 0.65595558277523, 
    -0.349481195125929, -0.274424055583514, 0.723475381322496, 
    2.12992700690101, 3.33042180284662, 3.88310800207882, 3.89661098003357, 
    4.12346597931558, 5.05096631182341, 6.59757158227971, 8.23105746249217, 
    9.22066214111983, 9.12504860264145, 7.79819580852841, 5.40137666217887, 
    2.58419882544332, 0.102439190730685, -1.68076532351325, 
    -2.63738431466293, -2.93041380106727, -2.68478538630297, 
    -2.02644936967022, -1.03291927355976, 0.310284336560999, 1.9771596736459, 
    3.50664912055247, 4.52713610022591, 5.01774881780674, 4.44879962943348, 
    3.10246105526469, 1.87876048189956, 1.35376240644283, 1.55650302880944, 
    2.12944538888888, 2.66823160984186, 2.91858215199028, 3.10620042402754, 
    3.51578207598799, 4.26801981442052, 5.3278787794728, 6.5212384560747, 
    7.63846349474472, 8.43015756683873, 8.63373558624529, 8.00280359066666, 
    6.52589188239452, 4.60639753834792, 2.58284050359336,
  -0.845077937413257, -0.00376754166089498, 0.575410583743149, 
    0.86202104606978, 0.881037611202352, 0.681042222902973, 
    0.300735555589698, -0.237739562912139, -0.861348086565226, 
    -1.43187483162843, -1.8426395910289, -2.1464590436694, -2.42109368003428, 
    -2.68674343897673, -2.97092090191843, -3.3053410034677, 
    -3.71339340622999, -4.1877719535434, -4.76593133310989, 
    -5.47432495527892, -6.26232543329271, -7.00031359227489, 
    -7.54715765110319, -7.79452685030905, -7.62890390714026, 
    -6.97347780555024, -5.95614276758121, -4.70340523022545, 
    -3.29012380118873, -1.91625749901876, -0.824877978606819, 
    -0.104040512726844, 0.237185025726013, 0.253532250896213, 
    -0.00686947291000328, -0.461827967408342, -1.03563011813219, 
    -1.65694196366043, -2.2732244746982, -2.81575162715308, 
    -3.18228986359622, -3.34991112868894, -3.43149900854854, 
    -3.53517364361908, -3.68408592979699, -3.87400934181103, 
    -4.12465883734671, -4.43995306801831, -4.79672941572169, 
    -5.19002816720559, -5.60868977774767, -5.99541847073993, 
    -6.23835324425841, -6.26706124535755, -6.0272106983023, 
    -5.47715603104317, -4.72729851197492, -3.88856684916465, 
    -2.92931329273249, -1.87084734982275 ;

 v =
  -0.112806168700575, -0.310410128353415, -0.559423157781429, 
    -0.849844272966729, -1.15336897179524, -1.43715313609338, 
    -1.66790068427652, -1.81349449726359, -1.83830533001875, 
    -1.71699126045535, -1.457136130368, -1.09511058116154, 
    -0.679757707683515, -0.258464508802848, 0.138695393052909, 
    0.495620678110905, 0.811369150436402, 1.09115046712602, 1.34880218677933, 
    1.60709411012794, 1.86922303625686, 2.10745771827726, 2.28303198949652, 
    2.36448433036527, 2.33781050616738, 2.18910474355979, 1.89893415771185, 
    1.4764575172717, 0.950114621550794, 0.351963278153529, 
    -0.260236646527293, -0.825069126666376, -1.3038850129587, 
    -1.66520907782983, -1.88009143900037, -1.93649122874658, 
    -1.83949639703967, -1.60552941290124, -1.26374830589903, 
    -0.86099544800694, -0.450584813838519, -0.0769224503495696, 
    0.224874821764528, 0.428213226999333, 0.522693892580878, 
    0.519673078782435, 0.452493983726666, 0.363221332016428, 
    0.283477842943634, 0.229753021161129, 0.205111203385768, 
    0.206754366317588, 0.227887301302383, 0.254177796436209, 
    0.27340568160676, 0.277900936909769, 0.260962208447883, 
    0.219406449231106, 0.147842260384438, 0.0387169934942612,
  0.744090375616198, 0.590163169054871, 0.289793796860106, 
    -0.202009434559132, -0.885906449634487, -1.68419429905407, 
    -2.46252606440557, -3.05806662458429, -3.34984655183068, 
    -3.2910885896123, -2.90028556000887, -2.25686892363625, 
    -1.49184827707835, -0.745310813227388, -0.121690788565541, 
    0.354046536286304, 0.707291379168297, 0.997829773847551, 
    1.29031963768244, 1.61584435333456, 1.99422261338948, 2.42458377766082, 
    2.84511031939474, 3.14607767113095, 3.23551465261265, 3.07292270436231, 
    2.66465265855914, 2.04949091871635, 1.29235810611357, 0.460071930390498, 
    -0.372449121671192, -1.10076485736056, -1.66458599765619, 
    -2.06828075714496, -2.3062403451665, -2.35183728736889, 
    -2.19143523515759, -1.83962747295825, -1.34950405512405, 
    -0.789946479006606, -0.220367487291614, 0.297715117510544, 
    0.69425787808315, 0.920187122430081, 0.964741440167793, 
    0.847559654124568, 0.609849366449775, 0.317347758377934, 
    0.0569953563455607, -0.105264196533844, -0.149096249089246, 
    -0.0886856685915078, 0.0433895333026149, 0.210120229721689, 
    0.373915731071679, 0.518251827149389, 0.629692786488842, 
    0.70532488466068, 0.762384980433689, 0.789098295641868,
  1.26270807697034, 1.17638382441497, 0.800582097768394, 0.0788417928036363, 
    -0.937455957556963, -2.10791676514085, -3.22933521088124, 
    -4.05934147781201, -4.41274518714007, -4.24977903685518, 
    -3.65209332712739, -2.71138770217155, -1.53575144502235, 
    -0.357604238540603, 0.555480851690828, 1.00449083850884, 
    0.984863961503917, 0.749987054499397, 0.669979728825767, 
    0.947063210748251, 1.5324604407221, 2.25620635395075, 2.91498354767915, 
    3.36347378110114, 3.52380320273106, 3.37293286729494, 2.88864362032753, 
    2.04110581057904, 0.978881797331435, 0.000573641484291296, 
    -0.744835479173809, -1.30805353138749, -1.71536416613023, 
    -1.96272082368766, -2.09344284959753, -2.09279573235646, 
    -1.88042403477724, -1.47467234609223, -0.956067370369909, 
    -0.336936123976876, 0.381877632992723, 1.09213736425504, 
    1.59689103730766, 1.70569134307912, 1.34378417839144, 0.666251679711876, 
    -0.0436792676778564, -0.596930336027946, -0.935950029979819, 
    -1.02267165152575, -0.837393303597595, -0.388948645454768, 
    0.187025722313395, 0.730464752801333, 1.09311280386712, 1.20695903895287, 
    1.16391255747923, 1.1075823307251, 1.11464608438104, 1.19281459980725,
  1.19657757677949, 1.14886475464706, 0.755168156178144, 0.0033475087451595, 
    -1.06109766769378, -2.26305461866838, -3.28301455929095, 
    -3.91028366832746, -4.11128028064353, -3.84987887583951, 
    -3.11388161249999, -1.96474112122563, -0.54301172260527, 
    0.738654302256832, 1.3626749444312, 1.23420012171969, 0.70189545375576, 
    0.208675495591196, 0.0807884762149248, 0.423434839349613, 
    1.26330863615915, 2.35799875879626, 3.29064647638321, 3.81252205033783, 
    3.90541432891427, 3.50358063080264, 2.56454292617386, 1.35731421793344, 
    0.135067400956721, -0.970988788629037, -1.74547182597712, 
    -1.98944309749741, -1.88569088494164, -1.76351386097118, 
    -1.72041704765791, -1.60179861085946, -1.30077843806164, 
    -0.908720275192401, -0.422551209588941, 0.259956567274765, 
    1.04178019263314, 1.61016999453272, 1.68849570914261, 1.2522898662034, 
    0.525392106307424, -0.254229826607117, -0.933995804385661, 
    -1.37310068770559, -1.42916354020032, -1.05779849887947, 
    -0.4625669156549, 0.203768786980536, 0.859399094937647, 1.38099599187599, 
    1.66581276616003, 1.58212251358034, 1.22715619304368, 0.933110740714037, 
    0.874550015350921, 1.0254328891779,
  1.0034855401937, 0.872258017705461, 0.433866624778387, -0.342260406914263, 
    -1.32491530889189, -2.22409280172987, -2.9061455217259, 
    -3.33139125513806, -3.42783461964895, -3.16436480302331, 
    -2.52456151570825, -1.48112489297782, -0.0870396704395119, 
    1.19256188516612, 1.67319720542465, 1.36756342542234, 0.716901471329893, 
    0.0800362894335941, -0.101120819446186, 0.42814468282074, 
    1.52606127902966, 2.78463447920157, 3.81749810454015, 4.35570905506868, 
    4.20779899892155, 3.37655195139007, 2.07940485914763, 0.437419049445323, 
    -1.18579421515411, -2.24692696711149, -2.65410996711905, 
    -2.42849639299503, -1.75378473935544, -1.12599913026538, 
    -0.827838206037851, -0.721591439238255, -0.685627510668456, 
    -0.59262995609705, -0.220840634549247, 0.431720410146386, 
    1.05374867013087, 1.31770359084619, 1.09378701450115, 0.45166050385726, 
    -0.392296813318714, -1.17536415604045, -1.67157159030805, 
    -1.76358474673211, -1.43740904187604, -0.832794423089487, 
    -0.113483906969961, 0.746831654157906, 1.64289944474515, 
    2.18999410401713, 2.0425037757389, 1.3930037384767, 0.807295864949583, 
    0.553249192532457, 0.616844410057165, 0.855602750036587,
  -0.0751930161917221, 0.104230235935447, 0.0161863144062146, 
    -0.45330042749536, -1.15402076826576, -1.87387053571187, 
    -2.43315701865334, -2.77479672693145, -2.84481593307731, 
    -2.63382359326875, -2.12302556059638, -1.2791821347993, 
    -0.153324730427887, 1.06493810903665, 1.9160138861201, 1.96690544275733, 
    1.24549875059426, 0.354639509857291, -0.0416693235952617, 
    0.252968321521278, 1.03280438481858, 2.17180930788562, 3.30673982537346, 
    3.89783920299902, 3.70520533184459, 2.79101906321569, 1.34080586397597, 
    -0.333420934676226, -1.66263772557163, -2.35912390230048, 
    -2.19445557917535, -1.21150272181119, -0.162789245445329, 
    0.209105106098054, -0.00794441892308186, -0.338065834441234, 
    -0.481218567271267, -0.388776551032594, -0.114914241516882, 
    0.254928818506419, 0.604080040322907, 0.780996733493252, 
    0.597484504260132, 0.0150608767013924, -0.821690020905069, 
    -1.67836292259554, -2.24380670054597, -2.23254081185161, 
    -1.54913909723054, -0.558176203068705, 0.286782325756681, 
    0.928569848799209, 1.49282992275196, 2.05444299862388, 2.24563043719198, 
    1.8607480601898, 1.25054725072164, 0.635890450083959, 0.0964978125296328, 
    -0.160664624926832,
  -0.770460232519185, -0.637815931866266, -0.444640862813761, 
    -0.501931349244252, -0.960383441307464, -1.61041976219418, 
    -2.05428052138862, -2.20379826101922, -2.16860964735358, 
    -1.95510953662876, -1.44915813945899, -0.634446004833096, 
    0.408839210496269, 1.27447933901431, 1.65033795016249, 1.85166089843325, 
    1.7777051948384, 1.23783171341009, 0.623504097274993, 0.306174690338435, 
    0.480466109364379, 1.21668871845295, 2.24097462619146, 3.00287447821972, 
    2.88599476299057, 1.66438413712663, -0.157575044732249, 
    -1.68409955256121, -2.26873203009891, -1.89550193439732, 
    -0.850812362381354, 0.101802765532672, 0.343857793086197, 
    -0.135909787887189, -0.773030420524463, -0.992472484795558, 
    -0.586141164213436, 0.0470665676316258, 0.459357590908919, 
    0.530064619853708, 0.378167480463121, 0.19753810399314, 
    0.0625790119253423, -0.156811747013062, -0.637773157290076, 
    -1.28551068149353, -1.76962543332252, -1.8451095913107, 
    -1.41577413680504, -0.538833534319764, 0.51171083123474, 
    1.27473604638684, 1.45844830351824, 1.24571058362735, 1.24938360764224, 
    1.61439956907193, 1.60795246232715, 0.930470010487539, 
    0.0301888941377847, -0.578467944672618,
  -1.04132769678598, -0.723981573687223, -0.214026233184181, 
    -0.138841884559351, -0.542237542064404, -1.19576169569251, 
    -1.70874734060296, -1.86329043873788, -1.76335763497888, 
    -1.4818357431282, -0.980405076174814, -0.249412102413639, 
    0.621902238608186, 1.48820100814847, 2.0578777104211, 2.06914965624641, 
    1.71288267182579, 1.28207449337462, 0.700846820625493, 0.220933910901956, 
    0.252884264650892, 0.77496910859096, 1.5331694962653, 2.16846390448496, 
    2.03845585726659, 0.677509429901421, -1.25389845278067, 
    -2.71341120286996, -3.05100356719509, -2.12024933541659, 
    -0.451771110214532, 0.715899111623137, 0.774082419431726, 
    0.0616199481144009, -0.666656354221658, -0.90492371322637, 
    -0.586469656945693, 0.0608563488032014, 0.639949075153608, 
    0.757601473175774, 0.44675596115658, 0.0405293321568024, 
    -0.127118321675491, -0.118328120421863, -0.32105238395654, 
    -0.747421971350311, -1.11999846971542, -1.15488628148497, 
    -0.669275876864775, 0.110125120732085, 0.843737862625193, 
    1.19898542834911, 1.15325747746964, 0.889046681594934, 0.550703447922872, 
    0.523103941100427, 0.718291010484214, 0.59456782526408, 
    0.00498238324653454, -0.698264267006351,
  -1.34431249269629, -0.67994053325066, 0.0184147130532058, 
    0.136364099642666, -0.300779427356113, -0.959760608659549, 
    -1.31561034921298, -1.32267893834125, -1.19429868256483, 
    -0.954744201280509, -0.654728496764302, -0.232349481449164, 
    0.433725217992299, 1.18113871289901, 1.77421660786037, 2.01337152925291, 
    1.67003037149909, 0.777608706650435, -0.181273383187314, 
    -0.759516371352515, -0.784809963311478, -0.0859554940207523, 
    1.07524533706599, 1.92677176759425, 1.52479514540865, 
    -0.00704193993243255, -1.53296205398716, -2.46685582930078, 
    -2.39459633310302, -1.2595858263714, 0.157324937858003, 
    0.923507267125418, 0.875766023654146, 0.325219440518089, 
    -0.187056029095943, -0.265269361217443, 0.140925117789274, 
    0.701074180423924, 0.878718850340112, 0.518859152204124, 
    0.00530787257824211, -0.281518206505361, -0.273701363755399, 
    -0.130613510444888, -0.186426204894961, -0.505590133052045, 
    -0.834463271582717, -0.828966009332418, -0.290656251662617, 
    0.578297558265078, 1.22593095252669, 1.18956555576475, 0.790369196934876, 
    0.533980112491692, 0.600175674088374, 0.856541414634842, 
    0.909617830592809, 0.401360058151673, -0.531543070100509, 
    -1.27948901721564,
  -1.3891373405309, -0.482666655494959, 0.175284413898402, 
    0.0891238067269797, -0.42771507294475, -0.918439532909505, 
    -1.01425292789597, -0.806013383068731, -0.556175563953308, 
    -0.405100603040445, -0.332269756887109, -0.153337663637758, 
    0.237142228026992, 0.837988997563358, 1.48883972637512, 1.83066245609459, 
    1.4913150292563, 0.279050246320348, -1.17991496005215, -1.95544128917431, 
    -1.72388517914609, -0.670814711865624, 0.73370209703046, 
    1.56948563060011, 0.921779431864895, -0.455295409703755, 
    -1.51843710129253, -1.8308295267798, -1.04998590421212, 
    0.233899001602472, 1.07023266829014, 1.06292164734733, 0.557493747046603, 
    -0.00709327458643656, -0.242310641492685, -0.0172191918409873, 
    0.577474932996819, 1.06614218563249, 0.882878358399315, 
    0.213133638710973, -0.38566638187018, -0.532990757359488, 
    -0.184186724607673, 0.0905074855000588, -0.18304713124195, 
    -0.680323737064832, -0.986143475374768, -0.782757836529297, 
    -0.0791487199744178, 0.782216493116072, 1.3011132543625, 
    1.09497025215741, 0.651085126053925, 0.48485534687145, 0.832949956760359, 
    1.50872967971862, 1.55136343302298, 0.502255814759141, 
    -0.809913625549158, -1.56644239485542,
  -1.02335997263915, -0.150022105476186, 0.226072857648658, 
    -0.0864893063234973, -0.654325102130772, -0.971093234710158, 
    -0.821959593194369, -0.462214643149215, -0.183376915675263, 
    -0.13179763389216, -0.228549676026687, -0.115023511801081, 
    0.335318964913771, 1.05622317179671, 1.76412311893336, 1.97476059254007, 
    1.10682785658252, -0.42778606720673, -1.66406305661173, 
    -2.14901459381941, -1.56141812660053, -0.289835305011787, 
    0.90753593561197, 1.19030319977802, 0.25306011127119, -0.814791755409963, 
    -1.37648411050647, -1.1858216175784, -0.074081710596973, 
    1.20101127163863, 1.6339542798533, 1.14673315629311, 0.412231554794374, 
    -0.194881672066088, -0.354674808791556, -0.0219071358036204, 
    0.562734142809992, 0.885247861051379, 0.523421875930554, 
    -0.147394048890554, -0.56748424507678, -0.503091945915021, 
    -0.0410656013028911, 0.12319413704059, -0.2856459018536, 
    -0.838127850825923, -1.11148601447572, -0.789803810858806, 
    -0.0345449694585538, 0.734463031108815, 1.00236526815433, 
    0.687620279146622, 0.353648971687119, 0.357678920099119, 
    0.969396045095236, 1.77358974384634, 1.57848741679246, 0.304428634738587, 
    -0.931853476944292, -1.44933709576628,
  -0.449917549782967, -0.0260455327292788, 0.00137142586337702, 
    -0.29940249497495, -0.746669976609888, -0.904718052720664, 
    -0.640620571002155, -0.274381656954842, -0.157281091250984, 
    -0.168862526070301, -0.0155739574872846, 0.422727326910126, 
    1.09941807354562, 1.69074073338759, 1.84189711804716, 1.36872029742428, 
    0.367357768733848, -0.613167598416946, -1.29636583511436, 
    -1.5014516032678, -0.873426050498239, 0.195330444290088, 
    0.76051769964738, 0.360530683263687, -0.457376456103888, 
    -0.910024308810281, -0.845002010125741, -0.349647052797304, 
    0.359443194079919, 1.02063651900746, 1.24362158084921, 0.89288354067894, 
    0.336407141526747, -0.0786625939150972, -0.204531385743167, 
    0.0234465158389805, 0.330573144241098, 0.195793538652825, 
    -0.24907304874615, -0.607404227817277, -0.65455572896473, 
    -0.408276704109344, -0.185348089202597, -0.13728920468451, 
    -0.24157738134481, -0.431203261853384, -0.464844193388143, 
    -0.206772258548924, 0.30209876255348, 0.692493001970691, 
    0.641610526328918, 0.411203767378545, 0.294225184519227, 
    0.445968530841749, 0.911200061477829, 1.14324399090566, 
    0.693652540174048, -0.162406575179783, -0.797163679432103, 
    -0.865315412528364,
  -0.151564922531556, -0.293127904502709, -0.451061351644897, 
    -0.54811021785242, -0.584174057653705, -0.443375369443852, 
    -0.128580253881297, 0.142482416084183, 0.0933355301653447, 
    0.0472666694016967, 0.38815799708926, 0.970694676944257, 
    1.35147807762025, 1.32067199022528, 0.817555838308121, 
    -0.0680102614578894, -0.662533195341458, -0.695207931872885, 
    -0.691222565396009, -0.68216305606961, -0.478056323498015, 
    -0.116610498142649, -0.0165792100181997, -0.402362187575008, 
    -0.640168167926735, -0.481556125547681, -0.185034279833722, 
    0.213205068018298, 0.574122491390107, 0.765138956928803, 
    0.812756697018083, 0.671522998360898, 0.350657857069886, 
    0.040784074055067, -0.114748304538706, -0.172097465140671, 
    -0.216354462105156, -0.384707464120369, -0.580925471607076, 
    -0.620661922875584, -0.597379396050287, -0.528084895867563, 
    -0.305700335843415, -0.0663910205231632, 0.0563054455934595, 
    0.172347560879005, 0.394091560262497, 0.610927195520682, 
    0.684021597198699, 0.568869792125045, 0.326227909794966, 
    0.224924270368211, 0.405817760027222, 0.653024910047661, 
    0.719121662209384, 0.43564122759614, 0.037239360775101, 
    -0.230432972171344, -0.314881733320055, -0.200930631846242,
  -0.212405783469453, -0.363929286003821, -0.497656703076499, 
    -0.579663964130946, -0.476127627294787, -0.17575882358247, 
    0.0996981026720046, 0.17660213109652, 0.318907687192718, 
    0.64134348804678, 0.808429907436529, 0.858383794568675, 0.7020307721444, 
    0.347215848376953, -0.139319896252857, -0.591035327848886, 
    -0.739199799903948, -0.681188340503093, -0.549731522475249, 
    -0.203970203579223, -0.0801522939244581, -0.414179699201104, 
    -0.662517815777843, -0.626374420125566, -0.382071948924842, 
    -0.105973377714493, 0.0543043084032026, 0.397159539814808, 
    0.818468626247604, 0.865558747367448, 0.697227494349795, 
    0.479186328273955, 0.181327178778995, -0.0852036043383836, 
    -0.242797725166852, -0.405420750081332, -0.533498503146686, 
    -0.554943759258196, -0.554042155677579, -0.537082596490502, 
    -0.402417183170115, -0.0664027276454464, 0.343310085291345, 
    0.535380707973209, 0.503377595886488, 0.4518914407137, 0.475100090423853, 
    0.548611633888787, 0.603345578495398, 0.574487429228777, 
    0.352661526246963, 0.179123727327497, 0.269676140138313, 
    0.370248362033569, 0.286100054109898, 0.0639816745045292, 
    -0.0797405823593192, -0.0637046851906198, -0.0516315845281578, 
    -0.119766115416835,
  -0.641628245504463, -0.4031997656382, -0.127232529343131, 
    -0.0499063669932976, 0.128490625573431, 0.392051868584711, 
    0.548623688697916, 0.822769770365547, 1.16919367004136, 1.18608028221236, 
    0.997490636882728, 0.917572788577796, 0.80644763088249, 
    0.604023039801861, 0.369890819133449, 0.186815811453425, 
    -0.106143390423496, -0.590331981352125, -0.825833287971561, 
    -0.645193731786593, -0.441352018948448, -0.518400560860782, 
    -0.591719023282194, -0.43480371117519, -0.273375153784522, 
    -0.189311322968118, -0.075628502938804, 0.126692892489703, 
    0.294784116597547, 0.342140367004528, 0.356361534746726, 
    0.297900409923321, 0.10607769821945, -0.142617669360883, 
    -0.378756465770115, -0.60715487575562, -0.765400020486381, 
    -0.729032849471697, -0.564256737466307, -0.439535513647428, 
    -0.266143382505502, 0.00882459520099774, 0.140983786201017, 
    0.0658667163905594, 0.00324801102570872, 0.0853316627749981, 
    0.203776707082338, 0.285165044262055, 0.400206772215657, 
    0.50613929506198, 0.465165576318934, 0.283934561327851, 
    0.062987950143452, -0.072106467164686, -0.0879115761979068, 
    -0.132341592852413, -0.241612974366385, -0.0889189071736704, 
    0.155407840578058, -0.23625430325268,
  -0.152901085499379, 0.15913126649865, 0.19105451069949, 
    -0.0256775341720264, -0.226346676676377, -0.412067803143106, 
    -0.662087234953765, -0.665846157036141, -0.256084959489332, 
    0.470538901925681, 1.09220018584464, 1.17277418434201, 0.943730277438035, 
    0.658912984449581, 0.354383926835895, 0.111644966403328, 
    -0.104352599114853, -0.3083923469162, -0.390625542146742, 
    -0.41327649170491, -0.380774566257086, -0.234924381876924, 
    -0.110703155821843, -0.0780540454218138, -0.164458124031082, 
    -0.284347896479858, -0.204895984165995, 0.0182480129720026, 
    0.29533696606457, 0.560147624748022, 0.653128882031376, 
    0.680461339294532, 0.633151572938453, 0.340612193797825, 
    -0.0763275443277414, -0.468884980995003, -0.779819770677443, 
    -0.905972488892877, -0.782729037393473, -0.476836102848239, 
    -0.179210019192174, -0.0811756178035447, -0.138553205571906, 
    -0.113054950190016, 0.113045661738804, 0.396352892715164, 
    0.592364909554057, 0.686240132358156, 0.574720747988766, 
    0.384801155760858, 0.45103617589229, 0.54252022923084, 0.308121469153075, 
    -0.0471830092634177, -0.277753930028334, -0.382547386737772, 
    -0.444296890763874, -0.424520409526698, -0.190797907211189, 
    -0.15537841615972,
  0.916646564880749, 0.803226437041146, 0.517092979124408, 0.269756229760973, 
    -0.152010129065377, -0.585308839047625, -0.625803451402566, 
    -0.37688597882698, -0.0997146034464907, 0.219233562857167, 
    0.505327062196757, 0.692085927349114, 0.709536068130787, 
    0.415209008702468, -0.0297009412037298, -0.361495996790997, 
    -0.437049736282296, -0.350669579982652, -0.376476268263922, 
    -0.501092747979761, -0.490241619591072, -0.249053217808117, 
    -0.0177979009675821, 0.00280791684907203, -0.169618105293287, 
    -0.412455022372021, -0.553716614086443, -0.456912431948157, 
    0.0389158480384089, 0.884038069556806, 1.54072131692727, 
    1.60047082356415, 1.1782051502611, 0.468032475279602, -0.208046119865502, 
    -0.6383590406834, -0.827386895175663, -0.775397370943742, 
    -0.528616033970037, -0.239985534565708, -0.0992895491700538, 
    -0.177030833201721, -0.380195249031741, -0.477237166001774, 
    -0.266988003036143, 0.0952464151757517, 0.361203755995763, 
    0.510983625680461, 0.555110271955337, 0.482383963339522, 
    0.400051441485056, 0.269441841022957, 0.0149213181788015, 
    -0.2768447167679, -0.447874298224482, -0.397467744615488, 
    -0.270519891891313, -0.323479268716717, -0.275922191823652, 
    0.386507066654798,
  0.541735048723257, 0.498779225163248, 0.574258801729002, 0.551564622617713, 
    0.125376317413001, -0.559930799618179, -0.992123024345792, 
    -0.781516650534638, -0.0967449209955964, 0.470266416892668, 
    0.61635899408723, 0.410032985754215, 0.154473739892841, 
    -0.0634861820677739, -0.292724759334853, -0.494232586754343, 
    -0.513104022347568, -0.345024645175564, -0.251385995318235, 
    -0.377221525345145, -0.595434655982524, -0.514332947151222, 
    -0.149068045471416, 0.175828643411916, 0.261294503401389, 
    0.083674879735868, -0.167281989978033, -0.258717996664532, 
    -0.0832657768492954, 0.418775661038186, 1.20705478040521, 
    1.82390480913467, 1.77424398396416, 0.962170168468766, 
    -0.133578491394419, -1.05462958782724, -1.55619144498217, 
    -1.41068985387106, -0.738252820566634, 0.0234239673409261, 
    0.461037350855539, 0.379659092488665, -0.0864570382116367, 
    -0.63013722120627, -0.97258171638335, -0.871549947012267, 
    -0.380963597429436, 0.165035518877336, 0.666542571576242, 
    0.982448298161112, 0.8947922031298, 0.493989791069885, 0.056077146074784, 
    -0.353777077241298, -0.60001402226994, -0.382811994733673, 
    0.102896839077713, 0.382686393893877, 0.372714662695419, 0.460001738988358,
  0.806295680677767, 0.677395641763558, 0.841554359242797, 0.890744781322697, 
    0.432058455797772, -0.551298403204489, -1.62876670832446, 
    -2.01720907215052, -1.21203841988236, 0.0260455232742489, 
    0.850559697223639, 0.702873818180277, -0.203202965187035, 
    -0.866941928468802, -0.811980177545637, -0.313602642105183, 
    0.0781227811117257, 0.166553827729358, 0.0355327255932696, 
    -0.206480908803457, -0.419239516157615, -0.392306934375581, 
    -0.118729554481426, 0.314029975655289, 0.565432175346009, 
    0.462627288697614, 0.16064975576281, -0.150772584223973, 
    -0.218101522942633, 0.108752092943229, 0.989930188735251, 
    2.01746343975015, 2.56556085855614, 2.155032970077, 0.654730080321769, 
    -1.23666165657104, -2.65292321510375, -2.88403469743095, 
    -1.89059032481605, -0.465098643806541, 0.636546430256797, 
    0.956905088725051, 0.401061638254664, -0.652411307801228, 
    -1.64483675883466, -1.95428617617995, -1.29500236626838, 
    -0.0816975730654661, 1.05543709214688, 1.68397596844006, 1.7567651723827, 
    1.29348085165756, 0.453728149802853, -0.365174731647061, 
    -0.954093390279899, -1.0670235236096, -0.538625645179082, 
    0.227226200092028, 0.897997303784751, 1.09081434637251,
  1.76452020474435, 1.83380944429894, 1.83784322024715, 1.55377857780926, 
    0.870525748879838, -0.417295852044505, -2.0309629479877, 
    -2.99526774184164, -2.30098558900992, -0.677208053696484, 
    0.584925159852826, 0.85602366789408, -0.142974450122128, 
    -1.47884273519203, -1.78081952843713, -0.989737458117681, 
    -0.0191843358783183, 0.541666766208999, 0.487347044136695, 
    0.0457626734188326, -0.429407472699388, -0.466797656363729, 
    -0.0209661898625792, 0.488912996094045, 0.547193655945641, 
    0.0215812287136694, -0.588860601155356, -0.865624775060251, 
    -0.722487952288911, -0.200983136235904, 0.878192229314402, 
    2.27112645045459, 3.16710677523701, 3.02517464753496, 1.68945326787805, 
    -0.449178087207767, -2.5048722872344, -3.28906919245632, 
    -2.41554430034582, -0.783935624005065, 0.587358134946291, 
    1.17524027606426, 0.744476274907502, -0.508557040326954, 
    -1.87605455324511, -2.51144021828589, -1.96058343443822, 
    -0.663072528005385, 0.749401270152291, 1.87858311589258, 
    2.39115343243319, 2.24133573607273, 1.48412561018376, 0.314222373589571, 
    -0.957767347758009, -1.81914882523245, -1.59103289189248, 
    -0.593162202482208, 0.547083518447271, 1.45971625755409,
  2.51778595061761, 2.6350162705495, 2.48802691883907, 1.99103046586357, 
    1.21031599334663, 0.0539531216283847, -1.49829877650728, 
    -2.70217511453629, -2.54123385024269, -1.25670166434536, 
    0.0376610473477505, 0.622391478811968, 0.0830851178049296, 
    -1.26713483336029, -2.2101605054746, -1.88060808877623, 
    -0.723594692441234, 0.395601887660918, 0.918079424623069, 
    0.741614136077861, 0.132704687811329, -0.160215029307497, 
    0.0242558641793635, 0.219106259192322, 0.211671208206164, 
    -0.327493600731893, -1.18196992420365, -1.61014252288755, 
    -1.36986798792108, -0.576064134141205, 0.596493090487595, 
    1.92110634688993, 2.89738165214303, 3.05290577433338, 2.23000517590887, 
    0.56721506230091, -1.33690854562831, -2.45819585181076, 
    -2.22190157108875, -0.997257639158455, 0.364836322560149, 
    1.12483039390945, 0.863191285393806, -0.292938384180741, 
    -1.7010307760622, -2.5299304992618, -2.30956487329914, -1.24909645559301, 
    0.130192468949902, 1.39618414088837, 2.21752854386836, 2.36056600239361, 
    1.7773903987672, 0.557696992465649, -1.02828195444997, -2.30755407200623, 
    -2.48018237552697, -1.33205152524264, 0.354550450109618, 1.80496211440398,
  2.20997332306862, 2.15170861144065, 1.93165251043367, 1.76565023518397, 
    1.36755526101408, 0.502797755808272, -0.681640234612965, 
    -1.66298512864795, -1.80488878975915, -1.05843769866499, 
    -0.0204186235584092, 0.649877069847489, 0.454741362056896, 
    -0.583910392005436, -1.64651901429419, -1.77475646503655, 
    -0.827617460997573, 0.512207368977401, 1.43544853866335, 
    1.53136544474902, 0.888019021840528, 0.182816535020521, 
    -0.160720178066613, -0.313555645466811, -0.43493256584158, 
    -0.79504680844191, -1.43338676117856, -1.88767265181455, 
    -1.76508911352454, -1.07933673756622, -0.0219758670398059, 
    1.27335945025608, 2.40865216866518, 2.83268884768191, 2.40731075568569, 
    1.39532115989887, 0.0850965941784374, -1.01238685841834, 
    -1.28836023233241, -0.58173943651713, 0.46037031942744, 1.09894505790225, 
    0.876392149434414, -0.207913370072059, -1.56766194433683, 
    -2.43594636977949, -2.49660050055059, -1.8388348859713, 
    -0.736398261756027, 0.377331616688498, 1.22861660315517, 1.6227714649042, 
    1.43351902344963, 0.618278564324813, -0.846125915924622, 
    -2.28135114549535, -2.71919750130685, -1.79521139845058, 
    -0.0835280209609241, 1.49427008011504,
  1.17737891329905, 1.62476183445604, 1.94138446690529, 1.91010159885397, 
    1.47165990049859, 0.969598321978574, 0.253961779836614, 
    -0.785041703124079, -1.24322560402477, -0.673307062406405, 
    0.240672572242823, 0.765282865416895, 0.567479211272455, 
    -0.313774436202449, -1.17929481064298, -1.23245981414825, 
    -0.433216079208447, 0.682395321783294, 1.51312999427203, 
    1.69651954588984, 1.12188371500597, 0.224269685122202, 
    -0.339846271121047, -0.541600587026114, -0.577516436395371, 
    -0.74936281595656, -1.29764467141401, -1.86697018093499, 
    -1.96864558967423, -1.44862559579733, -0.357613554553515, 
    1.03119565765316, 2.22014386339601, 2.8617657998529, 2.9080507877342, 
    2.29059702675213, 1.11715063758272, 0.11697719689826, -0.141289853476114, 
    0.284732910876511, 0.846131597536285, 0.921411457411363, 
    0.37438490451589, -0.51775830581609, -1.56545042548364, 
    -2.48233142839052, -2.88266160302564, -2.66066553936305, -1.769716599711, 
    -0.455445042434094, 0.69240665646578, 1.28754342887609, 1.20101546151269, 
    0.559082675362588, -0.500128009300358, -1.80587414898863, 
    -2.68120785987742, -2.40653040808287, -1.20213752288071, 0.229417318658391,
  1.54890249835952, 1.92745156062429, 1.8661097401729, 1.69152089443675, 
    1.2637124113936, 0.468054603786272, -0.297240476591724, 
    -0.66364436708522, -0.532741245557403, -0.0576990718991947, 
    0.383520379151122, 0.408519900097169, -0.112327041381919, 
    -0.834841204879238, -1.23588210538309, -1.01828620481523, 
    -0.268590559337342, 0.602383044055135, 1.12488058032337, 
    1.17798243224491, 0.888963056833356, 0.416425689062308, 
    0.0539902891495771, -0.210103703228092, -0.560713765275829, 
    -1.00954606191013, -1.45358290873526, -1.74458552542578, 
    -1.69899962216661, -1.16438465449234, -0.220131263336923, 
    0.834131066571907, 1.71906799362606, 2.21316598971294, 2.10800695062815, 
    1.47641367844971, 0.801765745372237, 0.537583551263382, 
    0.708075194324605, 1.01022554728329, 1.15646765452126, 0.919926804559292, 
    0.28389419323675, -0.743199468862732, -1.94754062762254, 
    -2.75589114563602, -2.86754130972587, -2.54370214500963, 
    -1.80489746454794, -0.58556422730582, 0.564017368106788, 
    1.24497311518632, 1.44891202182831, 1.17225700976871, 0.290152160277911, 
    -0.978973446510155, -1.99356116931678, -2.07040634312351, 
    -1.08770694326267, 0.38948212817154,
  1.78872498211226, 1.96489072767637, 1.56207309684324, 0.99518715954484, 
    0.406923034021154, -0.0842101667388026, -0.287699617808701, 
    -0.169346614944729, 0.0817473516483481, 0.232777289572203, 
    0.120049905767525, -0.249161154578099, -0.746937861993906, 
    -1.11491524948773, -1.07209548871021, -0.563374485116914, 
    0.195277638522895, 0.916251188425378, 1.43097877033278, 1.59283134854226, 
    1.39178142986257, 0.895953863282436, 0.152432838559445, 
    -0.60686964625115, -1.19660695417787, -1.64642193853048, 
    -1.93211311792481, -1.91593134980626, -1.5018120643127, 
    -0.779534968489438, 0.0674620923070696, 0.868732954743677, 
    1.31497717389839, 1.24389004729874, 0.992143749909647, 0.95760804470998, 
    1.12260762706476, 1.32696338730175, 1.55596623628396, 1.56672348575762, 
    1.24766883877097, 0.569858432890927, -0.463237683418743, 
    -1.5440850375107, -2.21284621186776, -2.29737845535709, 
    -1.89274834356785, -1.44627598467227, -1.39962407169518, 
    -1.20376580340975, -0.436781692404099, 0.406850941641686, 
    0.781190980938212, 0.590789476847938, 0.00485230477697449, 
    -0.645171975787635, -1.04674563315159, -0.986744238054595, 
    -0.306713145895125, 0.84240502795487,
  1.49439044863334, 1.59516661454014, 1.24302355834237, 0.669792953877425, 
    0.136845489867217, -0.18759565128532, -0.264813792940189, 
    -0.121361434638929, 0.15325033168884, 0.344881700045518, 
    0.206986957703513, -0.21355918065715, -0.586038984791002, 
    -0.636224370904096, -0.287444591124891, 0.364708217595791, 
    1.13547963608326, 1.7655862577583, 2.06715836861281, 2.02613920955731, 
    1.62520195982584, 0.867210131630763, -0.129071935490496, 
    -1.15135838110078, -2.00552414748331, -2.54358118705138, 
    -2.67340370065272, -2.41728726936307, -1.86630164997367, 
    -1.09741881458733, -0.268381870330506, 0.39687203273802, 
    0.814499733929327, 1.04020360848577, 1.19435169460923, 1.48473650796296, 
    1.99053868284766, 2.44145407715948, 2.64720844392954, 2.47934374667434, 
    1.7782450395496, 0.566426159106528, -0.752565375212689, 
    -1.68585425528905, -2.07341233864118, -2.06744427457647, 
    -1.88957604069024, -1.67678222763301, -1.49724337682193, 
    -1.30802904639078, -1.09240628246752, -0.852918799387949, 
    -0.616032888622469, -0.511467968018575, -0.56112353951944, 
    -0.658532403989383, -0.63874627886524, -0.332598376139355, 
    0.230204956225399, 0.941298619402047,
  1.13482621445975, 1.34713320259158, 1.17685919873216, 0.705276983269676, 
    0.18721966291995, -0.117922001596539, -0.152860394161338, 
    -0.0692555448871117, -0.00502822093401069, 0.044166393899835, 
    0.11170009459454, 0.17578332993988, 0.206451140103016, 0.25279536470904, 
    0.439389453624663, 0.849799882543076, 1.42846578037347, 1.98231738573237, 
    2.25382923372463, 2.08958396801688, 1.47500801016473, 0.541399009948588, 
    -0.499792737681012, -1.49534361134249, -2.34648116913384, 
    -2.9438327143777, -3.18325155135822, -3.01431283784043, 
    -2.47623710326696, -1.72155198308868, -0.942329278679277, 
    -0.249839166720374, 0.351211335598038, 0.871681687316174, 
    1.33477290074475, 1.83880509297476, 2.45073644034391, 3.03642352335592, 
    3.38136140347779, 3.32918345105452, 2.82969813463827, 2.01309601752753, 
    1.07048456066823, 0.101464137470333, -0.811655465012463, 
    -1.52651136247339, -1.93443622844715, -2.0557531928036, 
    -1.99704915333825, -1.89720815415426, -1.8200246565489, 
    -1.75169741400179, -1.6435796324095, -1.48047317511167, 
    -1.29486211864008, -1.07356085431322, -0.780867486733389, 
    -0.389675322047492, 0.0973576761239277, 0.650757694534632,
  0.439668508143221, 0.576201024913553, 0.585304587742149, 0.489510993760052, 
    0.337383030268616, 0.186644942739504, 0.0775003257356405, 
    0.0294211246964447, 0.0351750822314981, 0.0747786141267491, 
    0.144120278484629, 0.255336592028241, 0.435145877147756, 
    0.709245832835881, 1.07401316537466, 1.48383974949719, 1.85976505191147, 
    2.12037405331044, 2.17669221496065, 1.95768813185525, 1.46295122207425, 
    0.751884199868611, -0.0946686570489497, -0.97121349791284, 
    -1.76146760399061, -2.35925006672889, -2.69023368033943, 
    -2.73547679845003, -2.51881832448048, -2.07838887768385, 
    -1.46644835196778, -0.758160169446514, -0.0407497255209023, 
    0.634525697014693, 1.26651800793972, 1.85467424827876, 2.36532193370227, 
    2.74615306065617, 2.91668344875639, 2.81584802885615, 2.44410003404292, 
    1.86068847418966, 1.14946111873719, 0.420976896602851, 
    -0.212092738770886, -0.707653860882457, -1.08723785032613, 
    -1.38594784688983, -1.632582088937, -1.82031979375926, -1.93180829857995, 
    -1.98468023610066, -1.99449520008167, -1.94274507956255, 
    -1.78953703327793, -1.50820913440107, -1.11107078703183, 
    -0.650953163526828, -0.199298711316634, 0.176627365622219,
  -0.114451366447053, -0.0308021937798635, -0.00457259102196235, 
    -0.0216313030960233, -0.0580656505431449, -0.0915993870163411, 
    -0.104070675357646, -0.0829430802756144, -0.0244856348956226, 
    0.0698943988488687, 0.202571920339795, 0.383088925070767, 
    0.614744100205119, 0.884166877887425, 1.15988357009483, 1.4063097726381, 
    1.58856531729865, 1.67568931194417, 1.64074769896642, 1.4693408554753, 
    1.16179670210741, 0.734863210249909, 0.2258153873248, -0.309700373747217, 
    -0.806086080704919, -1.20589028716384, -1.47025385110462, 
    -1.57976941747714, -1.53311001871421, -1.34612444542263, 
    -1.04962428050127, -0.682844021875555, -0.277626047803656, 
    0.142030764825417, 0.552115966069059, 0.922916544231282, 
    1.22326958718644, 1.42704522540174, 1.51536070205431, 1.47551371298039, 
    1.30438878193667, 1.02168734019963, 0.673155665977384, 0.307003383180107, 
    -0.0459526615489157, -0.37007184915575, -0.649548503146215, 
    -0.868665331062824, -1.02109037743743, -1.11321194012854, 
    -1.16386969048573, -1.1843985262747, -1.17488075977319, 
    -1.12834234138563, -1.03923898969626, -0.916521207845838, 
    -0.771524010101255, -0.605975604821917, -0.426556449130036, 
    -0.253347128128928,
  -0.208352701465217, 0.196722767056692, 0.555058573379725, 
    0.823399010310252, 0.975139944527251, 0.994076291353205, 
    0.836317111711344, 0.494825606967882, 0.0454322315698141, 
    -0.424464446155893, -0.844666493171102, -1.16218785923988, 
    -1.33282422675701, -1.33552230245742, -1.16897999001694, 
    -0.843907440493962, -0.396726861258, 0.113612604438866, 
    0.675749069733888, 1.29549168478315, 1.9363994758614, 2.53140012245592, 
    3.01829250646623, 3.38379031683214, 3.59635725354547, 3.60924330463414, 
    3.39868828629563, 2.93044962058151, 2.18936425372244, 1.2460355780274, 
    0.166436369606712, -1.01508704414972, -2.20681872832462, 
    -3.29055834729045, -4.17926415089626, -4.79822516146719, 
    -5.08128744082147, -4.98209904538136, -4.49464585629602, 
    -3.65918979660113, -2.55153254747552, -1.29840236106303, 
    -0.0410687359231742, 1.10105183150812, 2.01031975300275, 2.5849584345729, 
    2.79181728882214, 2.66306632572183, 2.26087171768031, 1.65943998265216, 
    0.961050327767038, 0.265077093111754, -0.355176395336847, 
    -0.842719026693451, -1.17619165008266, -1.34055110486091, 
    -1.33534270800442, -1.18678048311455, -0.932368112694706, 
    -0.600417206623977,
  -2.86863554810202, -0.816434272603168, 1.48217785771627, 3.23389727984996, 
    3.8115117112028, 3.03150927585699, 1.2925746492893, -0.774779705426903, 
    -2.6246432720264, -3.76979024213225, -3.88130168929567, 
    -2.95466517409016, -1.35930335065848, 0.333059176072976, 
    1.58492781367326, 2.04211072083848, 1.70788350902427, 0.897750224602336, 
    0.00482745636276329, -0.446666933111156, 0.045464342135743, 
    1.62102427570844, 3.93162025252017, 6.20175735059234, 7.67882862485757, 
    7.93583344035787, 6.9251899441859, 5.07934589080814, 3.00706541916105, 
    1.05710758665643, -0.500816118969883, -1.45827250009517, 
    -1.99103504343542, -2.51438492899733, -3.32672181995128, 
    -4.50932541054422, -5.92649393137032, -7.26984425301513, 
    -8.10942569815432, -8.00735925177406, -6.69692597989505, 
    -4.16984075210028, -0.802810007003393, 2.67162488850916, 
    5.46796113541889, 6.9615369122963, 6.8109679502798, 5.16960935358841, 
    2.71695625923406, 0.375307667046957, -1.15768804624486, 
    -1.61620670126892, -1.18711808442047, -0.44570426238244, 
    -0.0567672298331666, -0.484495594314269, -1.69868650989034, 
    -3.14975972548548, -4.10984511216888, -4.0543008890194,
  0.872120228548316, 4.18902485132596, 6.15169915852172, 5.91615314218443, 
    3.88421800542448, 0.908557434265335, -2.64807933564145, 
    -6.37273933074414, -9.16225663493522, -10.0676053901698, 
    -8.88262896164561, -5.91988670578211, -1.65192435746999, 
    3.11170708825889, 6.72452829431064, 7.45263804361658, 4.60435321550784, 
    -0.238528263097417, -3.77227576137627, -4.00361205124688, 
    -1.65134765891405, 1.40952236268162, 4.10677843351019, 6.48711848802393, 
    8.60477679215771, 9.89208428924427, 9.41816518054316, 6.47657819990837, 
    2.06384969677265, -0.976181689587522, -1.24851466887855, 
    -0.0861922216126944, 0.820392108400278, 0.705423987608353, 
    -0.665795876328892, -3.19163288039899, -6.38537527545881, 
    -9.23052768069806, -10.5291324648327, -9.66294967293536, 
    -6.81430967124029, -2.67336774663964, 1.94733020126322, 6.13528005324274, 
    8.73694880519162, 8.71478004508111, 5.99176102031433, 1.56942916467512, 
    -3.03227247060181, -6.17929427603985, -6.59252202205623, -4.428311087882, 
    -1.19932504075274, 1.39526090932771, 2.46945638150372, 1.99124132801246, 
    0.398302990968048, -1.59935288920622, -2.79937245618951, -1.96955663330549,
  6.00576108437322, 8.78636703697096, 6.95793689836783, 5.8135647238338, 
    5.89342613967222, 2.53191406000636, -5.09857924388309, -12.2723383815675, 
    -14.2914286633277, -11.152101441, -8.01306111835616, -7.61085611566283, 
    -4.27916833994917, 5.81484208056439, 14.3024111952128, 11.8478566424009, 
    2.17154588885182, -5.26903800895371, -7.90939032065397, 
    -7.02367283812673, -3.12876911039824, 1.76845327543697, 4.43023373263302, 
    5.74127061216765, 9.16128226486534, 12.4615967229893, 10.4532654561587, 
    4.84871778230687, 1.56238909036379, 0.737903262973548, 
    0.0811203200308958, -0.0153132004510134, 0.417345270833948, 
    0.840452309957453, 0.964359309677833, -1.36804575013377, 
    -7.21621849061648, -11.8882148953004, -10.387278903708, 
    -5.55418757534905, -2.49595408972472, 0.373721627398358, 5.8465109702464, 
    10.0785774330486, 8.4795094118373, 3.23877652250225, -0.553351843203838, 
    -1.99447933548869, -3.84770845262074, -7.3287614380431, 
    -9.78501645731953, -8.02281618480268, -2.77233849919378, 
    1.81186095603451, 4.11670295593442, 5.47605321676573, 4.43217850860378, 
    -0.562879819229827, -4.31535532845873, -0.960054551520673,
  5.79536949773417, 8.99526894593344, 5.12429600261568, 4.69707777494285, 
    7.38757993542363, 2.91340731878193, -5.17936518078595, -9.10645124407379, 
    -10.8258187147774, -7.80501585613557, -4.18473855100572, 
    -10.0264166455172, -8.48101179129858, 8.58656213716803, 15.7846141626157, 
    9.41182635335235, 0.113635268161784, -8.56136773877882, 
    -12.0156069587772, -6.34218366826293, -2.04029690024933, 
    0.898626256216203, 3.86040431086884, 3.83181270878017, 6.92936781360763, 
    12.0482645000868, 9.46586421863353, 7.13676737465085, 5.2598529456177, 
    -4.65178256231104, -9.79090729968268, -4.50519435242549, 
    0.669293425390075, 2.5439174447626, 4.61498918376692, 3.55838316332809, 
    -3.73262560678954, -10.3681644157039, -8.13515300185306, 
    -0.86445923347433, 2.68489338266874, 3.76602444252424, 6.87428086446665, 
    7.68344668247412, 3.58028142380128, -1.69441943633296, -3.37208021853652, 
    -0.00921167671477954, -0.283561479230061, -6.91337367728482, 
    -10.0137366141114, -8.2877041111023, -1.79239625074889, 3.63184781420747, 
    4.03434654613919, 3.74548779538002, 1.65202421316053, -0.37039008596451, 
    -0.833254387522456, 0.0707552998513738,
  2.4383673889002, 6.14285610568363, 4.97062423637264, 3.31370427285941, 
    2.68751186096779, 2.52881982211468, -3.14067114618422, -4.69066460420687, 
    -5.46593130536149, -3.76709535804348, -1.89538929649468, 
    -7.76723704620617, -10.8766849083677, -0.613027491242222, 
    18.1227698885252, 7.92656306483197, -1.59788204047657, -11.6754347767406, 
    -10.9169345088711, -1.78251885112243, -2.5686888013415, 2.0671634105846, 
    3.87505851189424, 2.70041548823166, 4.25881534977283, 8.96529451415664, 
    9.89791908207816, 7.56856019259328, 0.636875449903048, -14.7868446248891, 
    -14.2074995230855, -6.79955315638444, 6.39492000332827, 7.2581993005178, 
    6.92092450588843, 5.90052441543824, -0.722810654366699, 
    -6.69449482549821, -5.94906633544859, -1.5280106482704, 3.32243831560822, 
    4.93643872136504, 5.99216652626897, 3.48202562025118, -2.02603387690835, 
    -4.6034771881806, -4.43075988909417, -0.848397531933511, 
    0.709401904128752, -0.519434114200977, -1.99959873559066, 
    -6.43307213530174, -4.31896435955907, 8.11194717005146, 7.39949664262313, 
    3.73535989704161, -1.16164203636736, -2.43252084638179, 
    -1.82603701226601, -1.19491086491449,
  -2.15011268207089, 1.07874956080516, 4.34015154011574, 3.24055690963597, 
    -0.727482635140738, 0.864473358249105, -0.323982447774227, 
    -1.86218066183877, -1.64094659193163, -2.3926997674978, 
    -2.80962917442907, -4.53911286106142, -1.99769523097228, 
    -6.22445453525034, 3.69256024933159, 10.916690942977, 5.53084267662702, 
    -5.11728037825837, -6.59178084938221, -3.62836261787262, 
    -6.85218870403784, -2.26209487618723, 4.3359340137411, 5.37724303309007, 
    4.67687733374652, 5.4378288815224, 4.34322001388577, 2.77441974892764, 
    -3.10793046738795, -7.44532618602625, -6.55637267448337, 
    -7.43992095594787, 3.25679840263053, 5.29463859972772, 2.3021024462516, 
    0.413435283613891, 0.266777211861836, 0.422874299491699, 
    -1.0915889995435, -3.03904286730692, -1.20716811107669, 1.99121028407146, 
    3.35305921147621, 1.5766515856644, -1.60154593464868, -3.03340913336031, 
    -3.79845316046044, -4.53459910728422, -4.98634389388868, 
    2.48034673550793, 5.2456429578531, 0.486531850693884, -3.74909424083613, 
    -0.197900674106575, 9.09041080868635, 7.60670275752646, 3.69943371677942, 
    -2.32519443726226, -5.3856191482824, -4.60822553611256,
  -9.06303444079172, -2.3399068462623, 5.69676799353043, 6.79722092778239, 
    0.349008837807131, -1.26766643432237, -3.17361689774699, 
    -1.50201169997378, 0.111452991285046, 0.179585195037258, 
    -3.20767620595936, -3.38873378609809, 0.906818542240091, 2.841414465734, 
    -3.27564146731866, 0.0861069407767088, 11.7928186029277, 
    7.69246553771065, -0.847088074752293, -4.14488850606794, 
    -6.1133941106139, -9.57066485689154, -1.77476479801227, 5.00497906460068, 
    7.7755440726704, 5.50146452784049, -2.12124420545643, -5.6096520764301, 
    -5.53009775855179, -1.89510927743073, 2.54110171305591, 2.05855417050957, 
    3.03290708023338, -0.562674810575073, -4.79492923873186, 
    -5.72181073431366, -3.34141422332977, 4.42518034873165, 5.66844684152885, 
    1.25084501520776, -2.20217398061755, -3.24966768118536, 
    0.594144395056994, 3.51211261313838, 2.36420104380135, 1.18545161407288, 
    -2.77945990605712, -4.95232500944092, -7.38064822581877, 
    -6.31763936037067, 4.7533173463668, 5.2864786058038, 0.978505533182822, 
    -5.40540469326745, -2.92191552635351, 6.51064818249477, 10.6220792784575, 
    3.71447376234098, -0.824247114189126, -6.64097005377523,
  -12.1396678647101, -5.20156696133998, 6.72650480491593, 13.4009717640183, 
    0.406568020711774, -4.68668701313217, -2.2922444634505, 
    -4.83129377602705, 1.85948780254525, 3.06700141126461, -4.67492115786333, 
    -0.601671842669539, -0.400099229150927, 4.06278968232848, 
    2.44603033503057, -5.5791036973934, 7.94099354481398, 11.0531958062842, 
    4.70767242293582, -2.301980942875, -8.54272446009535, -9.15210935307471, 
    -2.62957990976206, 7.18240631726994, 12.3303231708305, 8.25278844479378, 
    -5.523439197629, -16.4940036677155, -11.5850524497841, -1.69482251539691, 
    7.79038527547538, 12.7877542389846, 6.73833045845915, -3.57454121129184, 
    -7.92553780323374, -7.01187759720969, -4.50709794093985, 
    3.31946343001849, 8.71600705621887, 6.09094663253814, -0.749618858233165, 
    -6.80273855880591, -5.01391831714795, 3.88800609264078, 8.30412192372202, 
    4.28466424438816, -4.60429146240694, -7.28443253032176, 
    -4.12141101776943, -6.24899892544983, 2.44688777193655, 8.63814586626769, 
    1.01737988240071, -7.28061703010827, -10.2207704245458, 
    -0.725710277263295, 14.3079387115089, 13.4882304094984, 1.72866912323102, 
    -7.90625363842054,
  -11.4328044103967, -4.91459567097816, 8.21387963641582, 15.7570435497162, 
    -0.195435367216991, -6.4276974596698, -5.54662073422649, 
    -2.66936967421893, 4.04807879012046, 1.75602490303471, -2.43884359182509, 
    -2.22255550098886, 0.0374538152581133, -0.701704609896778, 
    2.44238150607815, 2.87315990782848, 5.1852892063921, 8.89896646048034, 
    5.21318014941062, -4.95364801471127, -12.5183604819383, 
    -10.4557130365398, 2.09310794019477, 16.0376240827488, 15.5925145563345, 
    7.58833432209836, -11.2709999305998, -22.396232068245, -14.2161237096458, 
    1.18867104734982, 13.7197439890053, 16.0927591594657, 7.97330521760559, 
    -1.05394012971676, -9.60744566651666, -9.30508761559407, 
    -1.53017221491911, 5.33959719107369, 12.3887367055069, 4.3168239936823, 
    -5.09612542659453, -8.43425643860039, -7.53013347944846, 
    6.76343681488348, 12.2458657923293, 5.11878073601294, -4.65252363422734, 
    -7.85460649587145, -3.88431325571135, -3.5594932124774, 3.51133486022999, 
    10.9229659054197, 0.0048292338098487, -13.5569632429105, 
    -10.0792110005482, -2.32946499566605, 17.5503198409983, 18.6404076827873, 
    0.908607963550926, -12.1825001596133,
  -9.37070324238806, 0.378460765037195, 11.0574085047262, 8.88522005053133, 
    0.156131862893055, -6.98970489668241, -6.12435884359561, 
    0.146805487315376, 2.93790289921163, 2.22470440207931, -3.56556012266636, 
    -4.82947538185715, -5.35275973542678, -0.251000650126093, 
    10.7484186781466, 6.36429347402848, 4.6150052748102, 7.56742395527653, 
    -6.85837329044299, -13.9269650977117, -8.56780673480704, 
    3.26308361898158, 10.4181665692975, 13.4600609027546, 12.6590529329204, 
    1.87807710827088, -17.7798147421334, -16.7219232137054, 
    -5.83748037087883, 4.77223305764667, 12.9886870954781, 15.7625997990682, 
    6.47141369331408, -4.94147973074598, -6.57314419482188, -10.963722676531, 
    0.0943175964007713, 12.3561483425693, 12.8850999704965, 
    0.449905609824053, -8.03244874823206, -11.7699985803093, 
    -0.417058181748977, 7.44880501174861, 9.59891985849706, 
    -0.347792219399445, -5.22208132660835, -2.42964341008, -5.0034746086922, 
    0.631220982185475, 5.89334987979066, 6.40668684971726, -1.96513354199096, 
    -15.8388565860698, -7.00942079334186, 7.87208004989888, 17.0010083778268, 
    15.4876622499429, -5.60534885286927, -12.2529366345405,
  0.201126156589438, 5.07842939367082, 8.66093577735207, 1.2127762719525, 
    -2.74524284029796, -3.51297963357452, -6.62240736610687, 
    1.73944916441598, 4.71911913893481, -3.12049920118967, -9.47984153137752, 
    2.310675444097, -2.42158259667473, 0.511324726853346, 14.4672540443776, 
    8.84897316234999, 8.39412273973476, -8.43152022230393, -11.4154621388119, 
    -1.33622578674676, 0.398017834826325, 7.54265991613202, 8.10725273279022, 
    12.0245166286451, 5.48838094610583, -9.27041267295417, -15.8319627816093, 
    -2.65202679627571, 4.98969011124907, 4.86760022075672, 5.87894768424084, 
    2.44720004135358, -3.69342985521006, -3.09335261490419, 2.99933112377424, 
    -6.12921925095719, 0.0360920754404465, 8.27414654752216, 
    10.4863911263931, -1.24964992374996, -9.31605452607572, 
    -3.67542960362273, 5.06193415632608, 4.30215359638836, -2.46361688553528, 
    -7.71268101902324, -4.88038471247383, 4.45634920770758, 
    -2.52035187796639, 2.61149414323087, 7.13171846155653, 0.51443603671788, 
    -7.2491550095065, -6.40285479324219, 1.76385654480366, 11.1767197319955, 
    10.4336118164032, 2.74056985215683, -9.7050678777699, -9.27173998458821,
  2.6210320826072, 7.98323864286439, 6.8865604510427, -2.2038959393453, 
    -4.44059370221295, -7.00060271399072, -3.86632919354759, 
    -1.61912433875526, 2.63028952448965, 0.207584431231517, 
    -7.82291263730603, 4.58990213601686, 2.36172091255653, 1.52434672985881, 
    15.4102960334222, 6.13717707081418, -3.99832734016118, -11.0825511922683, 
    -5.44140357366959, 3.0227603446381, 8.09926010392234, -1.03544215183223, 
    3.665937875631, 4.86644118074147, -2.86184772837697, -8.57428073428452, 
    -5.87100207479558, -0.934754474587884, 6.64341245360853, 
    3.02283826885254, 2.19358091464049, -2.17959151828671, -2.84485799128644, 
    1.14849256680801, 3.33789379679045, -0.109781000646056, 
    -0.514102483762854, -1.29432903251572, -0.322364124347768, 
    -3.28923623690086, 0.472341974875067, 1.86359691591579, 1.05001020233515, 
    1.79268027638844, -2.94309518826105, -4.34200235077701, -5.6345125345336, 
    -0.580301909699834, 0.90807194940299, 0.700361544033945, 
    2.21245398399647, 2.01726827981311, -5.489070208094, -3.83012006312309, 
    1.01035461488241, 7.06730453499819, 0.0369668328707986, 
    -2.61642219168899, -6.93415863062753, -3.43321423640459,
  2.46469058338119, 3.03878130115673, 6.84907718933897, -3.10449290311788, 
    2.40855867744736, -10.1869873107982, -6.16700271371261, 
    -0.241845140433821, -0.950181300740899, -2.16882728945048, 
    -1.43417151406445, 3.15103316930717, 6.15622741684483, 2.34999527599, 
    6.2442534946266, -0.630712741443872, -6.1805012288653, -1.91174975174332, 
    -1.67578705639029, -4.12760014636383, 10.4324011155486, 3.69201199050983, 
    2.45314764918055, -2.85439000738273, -4.71108312852081, 
    -3.32169209070724, -0.450501619905632, -1.30407195982606, 
    0.639476887191475, 2.11462544173952, 1.1876941162802, 1.73236449812189, 
    -0.280254964034064, -0.910976173977257, 0.571322837765649, 
    1.91310555691296, -0.249216716818317, 0.293775843778089, 
    -3.8480437672468, -1.72544029714287, 0.408233834628773, 
    -1.78129723951715, -2.21167683057674, -1.87164309448188, 
    0.00118584902383569, -0.944779169858303, -2.44384625910812, 
    -1.29694672820601, 0.0310389408996557, -1.34232327670931, 
    1.48727680278902, 2.56909078303031, -2.05449237166494, -2.79476656565539, 
    -2.6778451421286, 6.29955891015503, -3.60350868191728, 
    -0.380215400318859, -1.41495641998187, -5.22503845430495,
  1.61442537798597, 1.58462426470171, -0.494169345619772, 1.76741934345882, 
    -2.22627588899625, -9.28729885532215, -11.7468613304358, 
    -15.5110336852266, -6.63069730885739, -0.992704899514194, 
    -2.67350309146792, 0.0495404378992633, 0.866091979769105, 
    -0.630726359694402, -1.26367693028572, -3.71471698003134, 
    -2.91375235480764, 0.113184155459874, 4.51759433919648, 
    0.0423765124902258, 3.50563721641554, 3.32540004700591, 0.26832654837548, 
    -2.56575063819486, -5.89424207536502, 2.36906983740243, 2.70616845132429, 
    3.00045625806533, 3.65068434446823, 3.82348734484081, 4.23202838240843, 
    3.00440758125704, 2.07170643681696, 0.142761832859157, 
    -0.430216038806431, 1.56040787706372, 1.82014621218507, 3.09081531662377, 
    -0.55370927657593, -2.08775178768156, -1.2921603336869, 
    -3.61561077592369, -0.785671645462216, 2.18482113488107, 
    3.33557944534492, 1.67516675069387, -1.87719084727515, -0.44709281419338, 
    2.07892090790312, -0.375476668636416, 1.29665230044866, 
    0.793153668915268, -0.526866541497213, -1.52690745837257, 
    -2.86549135618171, 0.806612227358027, 2.17879323696587, 
    -0.803582755989905, -4.46479523709351, 0.793309351550529,
  -3.40506777298841, -1.3326466952465, 2.62937544573521, -0.465582541317677, 
    6.00754635178767, -0.529282948217369, -1.79857954064194, 
    6.30981808479149, 6.80827866792407, -7.05271534014783, -9.50537114938389, 
    -3.74625296322407, -1.22777032134393, -0.0875408811275384, 
    0.493927704499476, -3.30583263505503, -2.87253024887086, 
    -0.810426988845336, 1.41687481115852, 1.77913190079007, 
    -2.04020471913445, -3.24082287011834, 1.57642930551611, 
    0.537540100338409, -2.88468767349577, 3.2421229987391, 3.48524886847534, 
    2.64623011999202, -0.774383782146713, -2.34073750019726, 
    4.04568727977128, 2.77587958297553, 1.67312149407389, -0.975079850217471, 
    -3.02986354949769, 0.150858340953305, 2.81400124077204, 3.89097918806734, 
    2.42595320663109, -0.335924510136766, -2.77061572600902, 
    -1.52430578542951, 1.69406308477743, 2.80402115366015, -0.11182231418867, 
    -2.78314634695189, -3.30021381269724, -0.600294433462991, 
    2.17405932534822, 4.68844458325733, -0.619902186857308, 
    -1.77463162580772, -1.4310490781283, -0.243972710076943, 
    -2.07636861164881, 0.78026369679968, 0.61942358258975, 3.25586758248849, 
    1.8698094086854, -3.13688917654373,
  -5.71279400207339, 2.319061717375, 2.49751078467013, 0.901114063965675, 
    3.15606504637077, 2.88327462384961, -1.55324704833466, -4.32207404630619, 
    3.17001625545984, 2.36709561740029, -3.2685338533942, -6.58299442556724, 
    -4.29506338091694, 4.81078777478225, 4.53774996900867, 
    -0.681168283712201, -1.68399894175301, -1.69791402959886, 
    2.97797339524053, 2.38047560374801, -4.25648632154384, -4.51609844337685, 
    -0.775968580265268, 5.67093903567165, 4.40667150493195, 4.29193814117688, 
    3.22439367187842, 4.23041451658676, -4.93030199859238, -7.50149092384581, 
    -3.16657754798326, 4.67658833522426, 3.95838525832077, 0.890184959486529, 
    -3.34209307980155, -1.39157927799206, -0.745381885926307, 
    1.44972958297284, 1.55295176328946, 3.25928732495335, 1.61389652677237, 
    1.28811390694278, 4.35193875264289, 2.5257922505563, -5.80709750101094, 
    -6.0009680088838, -1.1900381763361, 2.6232181062824, 6.61761993187276, 
    5.27381100292101, -1.92498361666748, -1.61239283122538, 
    0.135652767027902, 1.10492764969509, 1.58880809847199, 1.16334367413839, 
    0.909826871247745, 1.60239946743608, 4.27509114985907, -13.04626783172,
  -0.64123206972958, -1.16620132992775, 0.971449569383866, 0.977875733684621, 
    2.39732137687908, 4.81708529868364, -2.45653194381107, -6.89621028409993, 
    -7.78462164130571, -1.07286885619625, 9.40928407787643, 
    0.762462633576023, -7.0175937570319, 0.0190607288201972, 
    6.27796996969257, 4.15820637956452, 0.0176593248328684, -4.5041873763327, 
    -0.449665877011881, 4.47470376752275, 0.175638345025305, 
    -5.82209797676616, -4.9723011763148, 5.12422695824113, 7.30828119756198, 
    5.63149140414143, -0.943973298912371, -1.85355693114813, 
    -1.80164268659693, -7.09949684603722, -7.37735383338399, 
    0.863312613807102, 13.1066135516859, 7.91929695186669, -1.93587024554416, 
    0.34969086411649, -3.2524063700336, -8.4676086315774, -6.3113279005812, 
    1.41869097574463, 6.86764970444492, 7.10081536814529, 5.50983205809335, 
    1.4433496678523, -6.00491119747633, -8.30901532814025, -4.57194687558314, 
    5.79539335102322, 6.67416549481584, 1.27666793493501, 0.799123273507739, 
    -1.0731369701883, -2.02323048843125, 0.80948800144633, 1.39436635546725, 
    2.0082044000702, -4.2229209493477, -0.531718309286015, 11.0605255992291, 
    -9.96440625007372,
  3.11152371193222, -2.22108463106588, -6.34371118869362, 3.98414261701737, 
    6.7973537984621, 2.4390149074321, 0.281650887158671, -11.2958489555319, 
    -15.4425630199142, -6.46920790250436, 11.7235989812043, 12.1222825726585, 
    -0.826784894072352, -6.48977824668707, -1.91467386203842, 
    3.22080065058096, 2.48630581056855, -1.89293189658966, -3.73106670171515, 
    5.87770706015275, 2.95079527453217, -6.693056744309, -5.79769287692377, 
    6.34076636356755, 5.36273409683732, 1.79730382723216, -1.07081044752609, 
    -3.03402637751851, -4.65310212065372, -7.08283591339332, 
    -2.30235367316474, -3.94253418162219, 13.218141944999, 16.2705010054209, 
    6.46631242902744, 3.85932122448237, -7.22354395248746, -18.5773227974568, 
    -16.4405964384951, -5.7636172344957, 10.7825799848769, 15.8631566688872, 
    7.32772185319259, -1.69799410465878, -4.72512034048733, 
    -6.54544323027933, -10.8275311413566, 0.157509040154551, 
    6.41092722241014, 0.775884743217355, 5.43407295601693, 5.39242581474342, 
    1.53370672549412, 1.6745555838389, -0.247952898296459, -11.3290171173983, 
    -11.7950951631278, -3.86615242206208, 11.5233320119596, 5.12872699559541,
  5.0766092074388, -0.380182027089983, -6.14257307544852, 3.32267001071753, 
    12.9773417859493, 9.4811065206037, 2.10320787932814, -14.1674786192045, 
    -21.8034334938984, -12.3918618723941, 6.39648329003926, 18.7136578372625, 
    11.25433759427, -1.85247839945924, -11.8222192629854, -12.2082760582605, 
    -2.9293842052485, 4.95330943991486, 4.96032073608054, 8.92637722945231, 
    -1.3966687471154, -9.62137927806673, -9.14770775686048, 5.94171098654199, 
    10.1162110167977, -1.8788069480514, -2.34425561907668, -4.2531627231856, 
    -3.71752724034655, -3.24183923594111, -5.39750833335371, 
    -3.92496923994237, 5.0652937955661, 17.0520166494368, 19.5226944876023, 
    9.71300200699924, -5.86820412193382, -21.7371171464002, 
    -21.0907487121257, -8.3944848179436, 7.18262949943723, 13.4403361759214, 
    12.3741315713404, 4.19424011685419, -2.38451887371071, -6.41070643055622, 
    -12.3842287502057, -10.783005200052, 4.0081786307306, 5.0585149165957, 
    1.50635775504664, 7.94965361975654, 9.11792287727593, 3.19894765476748, 
    -2.57026406270742, -12.2599928577112, -13.6476628849474, 
    -8.08459109007048, 5.33432441518901, 12.5779396435234,
  4.57448483573027, -1.44344713194911, -1.27868365449711, 1.95763693326236, 
    12.2391950929776, 11.4505941373661, 3.05230915040451, -12.5011017196397, 
    -20.2198458329727, -12.4347137509981, 4.93065544064075, 19.3935337685808, 
    14.957079013614, 3.43565398482262, -14.5199393649622, -18.4196021764341, 
    -7.71172223771052, 4.75614177602356, 9.96170218041402, 6.44838395737773, 
    1.65515539385944, -7.82507308460977, -12.2470702965797, 
    0.724685949310121, 5.73304671297477, 6.50395247182054, 
    -0.378675483651902, -5.44484808183494, -2.99239180709513, 
    -3.04406398072178, -5.46619769844312, -4.49237882783702, 
    1.11142247440391, 12.1108350441047, 16.1108823265278, 11.7262212945818, 
    -1.31039548196239, -19.0864794181518, -18.5049016283071, 
    -6.90046470463585, 4.39538355093625, 10.0367408121306, 11.1506051745508, 
    6.51356704102606, 1.24354160242521, -10.1458325945725, -12.1524532614452, 
    -7.68712862392665, -0.423171598303786, 1.27150826994484, 
    3.41429844563042, 3.28961723914112, 7.82665243003923, 6.30464748979045, 
    -2.2665584665733, -6.1023558109798, -11.1475750490686, -6.70252054772397, 
    2.30925462685332, 8.37797466829942,
  -0.870193721950049, 4.26003536910225, 1.22530692714337, 1.18634869284561, 
    7.84631106827774, 10.0252856592775, 4.51853545880897, -9.30349959809719, 
    -13.3497014572639, -6.69092719187626, 5.75522818042558, 15.5646619592022, 
    11.2253283476569, 0.632850230032405, -10.1349785894114, 
    -14.4428634696905, -6.73763414392273, 2.70051729398472, 6.44992647341278, 
    6.94682071892971, 2.10278407294184, -7.99071644520566, -7.97047471900776, 
    -1.67437793637233, 5.2449089952321, 12.2418349389912, 0.104264567987852, 
    -4.18405271733718, -4.53406384247528, -7.06658853745738, 
    -5.49475371349166, -1.68197659644397, 1.19021940779452, 8.20017140032624, 
    12.660603115065, 11.8831519546865, -2.01048199156375, -14.7410256215491, 
    -10.8158399271289, -1.71486994266406, 3.71115006689687, 6.37022208703598, 
    7.18780176396607, 7.50180542258753, 0.119996989448852, -10.4689220610806, 
    -11.8300881700858, -7.36716569964636, -3.27909534957293, 
    -1.58568072634052, 1.52196141095844, 2.32253678482361, 5.57240267844289, 
    8.77206573293975, 4.38841572728836, 0.567518749299361, -5.83073555180863, 
    -10.807351615366, -2.32666950929227, -1.05605328433436,
  4.19826091502177, 7.17178111822106, 1.55376435022423, 2.02555487255696, 
    5.0811453148433, 6.2689188647072, -3.20801482982044, -8.97327018734661, 
    -3.20300532675963, 0.978670091007765, 6.62971717017783, 8.33108242183598, 
    3.91607385677027, -3.76133749397614, -7.24678877322924, 
    -7.66188185851958, -4.12342914132459, 2.17439853071502, 3.70700065816561, 
    3.41085962980887, -3.51725156566088, -0.678861415196236, 
    2.54196779402709, -0.86514928838048, 8.21312158188901, 6.39289969391542, 
    -0.845004757722787, -2.53311384613101, -8.27939241369507, 
    -4.69008791783318, -1.97185712154822, -0.246485819689939, 
    2.84501120191432, 6.88797274937659, 6.89297660437203, 0.804347250612281, 
    -6.3348360863901, -7.95945548825247, -0.942484497236776, 
    4.63111315259145, 4.95618304621172, 4.43187094298268, 5.98227231077334, 
    4.98596558042293, -5.04757925814985, -10.0095078364661, 
    -9.66069830535562, -3.66509281347351, 0.0676618909750648, 
    -4.12160634236036, 2.12146613510891, 1.7430372960314, 3.81808223948091, 
    9.34826230784225, 10.8200837603232, 2.03507150072304, -8.97471330095299, 
    -12.0787277216986, -6.31691179624518, -2.398652796974,
  13.4913393819634, 3.8715745703998, -2.74419331721599, 0.675713767239428, 
    1.8940375945794, -3.18036173862003, -7.95642586613488, -1.67261601364155, 
    5.2750004822005, 4.03368871934403, 3.94300383889419, 2.19623664268074, 
    -2.56616980733188, -5.39361741246023, -6.85580069794476, 
    -6.65000501357339, -3.61564439424354, 2.6631478061962, 7.07332996760064, 
    1.19294707144712, -1.73279607915946, 8.27760503637534, 7.74400093765536, 
    0.52353766333543, 0.829581911073558, -1.55742456979299, 
    -1.04592623722163, -3.65639848124117, -5.3415377321401, 
    -0.615823468809279, 2.16409397643516, 3.73802852743421, 3.26424585576829, 
    -0.600741691585757, -3.37658111413231, -5.59566322733752, 
    -6.43833125596225, -3.25575031843086, 2.86290604131225, 8.96393275218473, 
    8.36303304960853, 7.51418777964686, 4.01701626194896, -4.01493984169087, 
    -7.15236312483182, -4.43832924167011, -0.274962923760025, 
    5.93096023155292, -0.194930718647427, -10.0222955607334, 
    0.599088638181558, 2.69535898800966, 3.90217568660146, 4.53284003519595, 
    2.17071420901432, 0.00867417155601753, -4.40485210970439, 
    -7.49395419193502, -5.09290818148417, 0.991129383276749,
  10.9117207149762, 5.31681828590112, -2.85729000160844, -2.17400109729018, 
    -1.55019780532191, -3.79841704228287, -4.3586184484863, 
    -0.714189928177273, 5.18313290881012, 5.901337178126, 2.28352893848091, 
    -1.46050096259512, -4.14619810086888, -6.0655779950703, 
    -6.67637843554884, -5.96516724378686, -3.21424860229879, 
    3.37359650484698, 8.43423070406056, 7.40365008755992, 7.41114591660111, 
    6.18209001448092, 0.322336781184128, -2.12034712385481, 
    -1.68716668750921, -2.35221467999242, -3.88740858199969, 
    -5.32020990833578, -4.01742657577689, -1.16682969921383, 
    2.30559161370606, 5.38148196485807, 1.74673753958932, -3.468885129694, 
    -3.60424796395058, -5.01821828846907, -5.28396404484205, 
    0.29498078280255, 5.80849306940562, 12.7192143247833, 14.3265588501572, 
    6.45999591607124, -0.845991118446604, -4.41580310954898, 
    -5.6323551219511, -3.48383355134491, 2.39351870898801, 5.03765529506317, 
    -3.02248136823511, -9.27596011953388, -5.77519143071811, 
    -1.30109127173291, -0.866751776846689, -1.00906811105732, 
    0.113842019379674, 0.832867197823508, -0.502292903927766, 
    -2.74070200514338, -2.63075416223822, 3.39360405738388,
  7.9475757411792, 6.03712292946055, 2.17116752451729, -0.758506280488752, 
    -3.05831797554426, -5.88890494313929, -6.70763320480755, 
    -2.84734720112264, 3.15823405794875, 6.2031415444481, 4.78470309576616, 
    1.43181170801746, -1.61088755038892, -3.68023123701237, 
    -4.23511219309382, -2.64862017214239, 0.619055539093065, 
    4.47217884471065, 7.50169719023837, 8.18389238988001, 6.19206954647904, 
    2.93387252156909, 0.744619130751379, -0.0122228265205423, 
    -1.21607679484206, -3.97753031351196, -6.98111758521192, 
    -8.28746665753086, -7.26896713441111, -4.71395203067795, 
    -2.22526079230627, -0.700105694082884, 0.596416975872058, 
    1.71769622668444, 0.608782132640827, -2.15118236674778, 
    -1.33022471350475, 4.88240365224832, 11.6203519880689, 15.2000299503871, 
    14.5987383827119, 9.09004358982505, 2.4105636408123, -2.28926421055547, 
    -6.38301337298805, -9.590080990125, -8.5192819199367, -3.33821189273007, 
    -0.0347977807462561, -2.78902370762008, -7.37144636357133, 
    -7.33846878176317, -3.81691444694367, -1.18143296881599, 
    -0.755338391940308, -1.86401931367975, -3.19446296141759, 
    -2.59461116997745, 1.08412925775156, 5.74111045797702,
  4.74733062249814, 5.79775749200435, 4.73875494833793, 2.05336648248866, 
    -1.44968597035731, -4.54464072028819, -5.93522032704959, 
    -4.85899377770829, -1.59228337835672, 2.30572155016921, 4.80242316030423, 
    4.65608098793328, 2.33335497994895, -0.0660704362909539, 
    -0.326267791633297, 1.99626912636188, 5.25538005406784, 7.40659464513863, 
    7.89134629838733, 7.1815863307984, 5.94001145271861, 4.63921351517291, 
    3.33742497894816, 1.61203273513635, -1.14259836729417, -4.92179176367598, 
    -8.73284092542272, -11.1997081156904, -11.5459873634695, 
    -9.94946632557868, -7.02565574167441, -3.26550860169291, 
    0.559667672146906, 3.11265884521945, 3.41098198254373, 2.18252031386632, 
    1.60001228561529, 3.65721026884853, 8.11783581216372, 11.9604644862581, 
    12.4158185821428, 9.22148698742346, 4.07418981926568, -0.946833494061982, 
    -4.62072693350415, -6.72670117337932, -7.49353444091909, 
    -6.9133071624652, -5.11116182462652, -2.89649779846006, 
    -1.28475160385264, -0.918723720612281, -1.52553476605565, 
    -2.568702196337, -3.89956209171564, -5.24921032956394, -5.8214251019129, 
    -4.79808143432023, -1.96520660591634, 1.76800113896212,
  -0.426640178456187, 1.42929441739459, 2.23527666902231, 1.82971551209949, 
    0.520719882715169, -1.08307553645803, -2.24343563062539, 
    -2.3887631527164, -1.44865864175496, 0.126706129941063, 1.6079524605546, 
    2.44899534680692, 2.6177306865615, 2.54441736761481, 2.8092256080657, 
    3.77954693553842, 5.42173078045756, 7.26186700834411, 8.60305083280447, 
    8.9415263207221, 8.12732620438763, 6.29961964600271, 3.73292603021306, 
    0.721487407568701, -2.4463762024458, -5.51016456103297, 
    -8.16868142568135, -10.0402261386796, -10.7571518469109, 
    -10.029949700366, -7.80957737931927, -4.5685780955448, -1.19885796320628, 
    1.40079789765165, 2.74741977586283, 2.95416133778769, 2.61786832205616, 
    2.38252344067868, 2.62573831523304, 3.36231293247422, 4.13121330397915, 
    4.25165731252875, 3.35145242321592, 1.6130124919303, -0.349352229700211, 
    -1.87899926116438, -2.56388114736031, -2.31820825741304, 
    -1.32542108044428, -0.00650422196941631, 1.09132071128186, 
    1.48995384516845, 0.812152009877541, -0.929223552131446, 
    -3.19774939267349, -5.24341933138702, -6.4145327553724, 
    -6.31005748613099, -4.96052107843093, -2.78899882004564,
  -1.76782502306405, -1.30383072491746, -0.822260612179789, 
    -0.369762868778222, 0.0238057746636031, 0.364870287510031, 
    0.658264735007648, 0.895670162010119, 1.08509815811335, 1.2502478216856, 
    1.43277793112593, 1.66405939450713, 1.94852350101581, 2.27024515207866, 
    2.60796962112701, 2.93479337580967, 3.21940950814606, 3.42061672590735, 
    3.48820597614837, 3.35793789022659, 2.96940877239738, 2.28645371416095, 
    1.32079974641837, 0.128671953346047, -1.19232586950071, 
    -2.50588488805601, -3.67493337155199, -4.57053181213083, 
    -5.07552952609372, -5.14088830423576, -4.80506473821033, 
    -4.13475445321241, -3.20665171146805, -2.1187191054236, 
    -0.986434769078468, 0.0891653076472836, 1.02493185484467, 
    1.76713151577718, 2.30526391033857, 2.6399027170323, 2.77634550817349, 
    2.75088298728291, 2.6083859391238, 2.37155474987563, 2.04094009171492, 
    1.63093025998324, 1.17795170895515, 0.722265067035203, 0.281170035416676, 
    -0.141845660503047, -0.555470636560469, -0.987182743820395, 
    -1.41206984192665, -1.79161167841589, -2.11374618174595, 
    -2.35530355392951, -2.494426521529, -2.52670881970976, -2.42193427189264, 
    -2.15876746453339,
  -1.46451220622127, -1.64119593143673, -1.71355956964674, -1.68433294404149, 
    -1.55974090540727, -1.34553246860248, -1.0900640653484, 
    -0.857588294242198, -0.667028745119074, -0.52206975101005, 
    -0.424526111420916, -0.370106797978641, -0.338152701284067, 
    -0.306792305918805, -0.244302280341491, -0.111232033761018, 
    0.111132627826909, 0.404519739139451, 0.759752227862249, 
    1.17437189160878, 1.61629508239294, 2.01958383388544, 2.31772620746334, 
    2.48884860178333, 2.5178118896464, 2.39448685381834, 2.133857980417, 
    1.75852361757622, 1.27136520120823, 0.72546586842622, 0.184524510635378, 
    -0.345753979072765, -0.847418611245744, -1.28393874380207, 
    -1.64899652279019, -1.95361666004443, -2.20517968480707, 
    -2.39283130002455, -2.49756549087232, -2.49228495217133, 
    -2.33592539915312, -2.02291000377854, -1.58423838206919, 
    -1.04050240282617, -0.415196085867543, 0.228516905395331, 
    0.824477342552581, 1.33503263329354, 1.73398864573296, 1.98775534516121, 
    2.08168245944792, 2.01777224764493, 1.81121946214353, 1.48974906562256, 
    1.07697691134314, 0.612607209457531, 0.130613870395259, 
    -0.344567721516718, -0.789596234954549, -1.1759156406916,
  -4.98979259298961, -3.88088671749721, -2.01476680643861, 
    0.0778577467148643, 1.75061025056363, 2.50445156147738, 2.26068572372177, 
    1.24515513506654, -0.238755336199873, -1.72124267449366, 
    -2.64309607992202, -2.64348402709274, -1.78320136865058, 
    -0.456882386498475, 0.797556297981761, 1.5240009917776, 1.57518462276583, 
    1.15057744986803, 0.490255751592384, 0.0151946892539194, 
    0.251340415197312, 1.45204342971047, 3.43345399059882, 5.55091157780396, 
    6.98956902314726, 7.14423290440683, 5.89319819219244, 3.69097197543709, 
    1.4130182498706, -0.223892541374413, -0.907870068684978, 
    -0.643929199288822, 0.162002592565032, 0.827139601727904, 
    0.744825308167045, -0.383747692219864, -2.46939361821846, 
    -5.08111124423155, -7.52013820524522, -9.01828863635611, 
    -9.06902182524004, -7.53051602241585, -4.64946146314484, 
    -1.06308224832791, 2.45251789737273, 5.241430927695, 6.78120785941526, 
    6.79974390151717, 5.49721765851421, 3.53254637602669, 1.66578402224402, 
    0.434360911837921, -0.0319187599706038, -0.0158686481260515, 
    -0.0125917159103344, -0.497453996952456, -1.60209143157551, 
    -3.06034088364934, -4.39774447757121, -5.13805862880598,
  -1.12045761266858, 2.13087277967325, 3.98259821176242, 4.34720599522312, 
    4.17507744816384, 3.71825832406019, 1.95764259108954, -1.64891683601292, 
    -5.60776129746767, -7.9656716008687, -8.09903273527092, 
    -6.54177965773418, -3.69120498980394, 0.283763766228013, 
    4.45781464639654, 6.82577238272445, 5.77125049991326, 1.72639757572482, 
    -2.29294510524181, -3.57771839426712, -2.18860085200469, 
    0.12668698559167, 2.38327467788392, 4.83476828275948, 7.44548298278942, 
    9.08155854912015, 8.36391382764423, 5.1042174963431, 0.782881742314945, 
    -1.94037995368375, -1.52212233554929, 0.894761940237196, 3.352916496202, 
    4.67914433891572, 4.06218425235988, 1.00137659350255, -4.07443979337658, 
    -9.37954683782871, -12.5852657676349, -12.6656682829248, 
    -10.2988221571308, -6.58377554532019, -2.03575458008294, 
    3.00129206856087, 7.42134361662092, 9.38231741563201, 7.96572229823045, 
    4.15617820143505, -0.193132086515186, -3.47745700537521, 
    -4.65017910377492, -3.59576351959113, -1.20132508338998, 
    1.11273685825218, 2.14005813047156, 1.42452082058035, -0.676098267341479, 
    -3.23689451972839, -4.81709803289088, -4.04704888245937,
  4.89773762350929, 9.39007889015408, 6.38981555800446, 4.56229285368312, 
    7.51453735663693, 7.34958549842352, -0.331881933319451, 
    -8.43883457129875, -10.449485574226, -8.88181883338837, 
    -9.08777957386695, -10.9127927743062, -8.53315655039986, 
    1.28623997514466, 12.1952229588542, 14.4491813137239, 6.38113756688471, 
    -3.50550360634266, -8.63457918109456, -8.76482082089544, 
    -5.43790279612321, -1.0427332613402, 1.46220941401288, 3.04943686333854, 
    7.478578941118, 11.9883773574613, 9.99799795567857, 3.6208807953011, 
    0.896634114164186, 1.98533707849049, 2.12770058174841, 1.50711251223425, 
    1.61455818372543, 2.39982866961433, 3.27468454920952, 0.978800664385147, 
    -6.72061499166007, -13.6475416306942, -12.7873618786239, 
    -7.99285649973035, -6.073180092033, -4.1703837786994, 2.78018090899446, 
    10.1816434911321, 10.6715383093376, 5.5538431461722, 1.43156960250058, 
    0.529329917538082, -0.700276713424433, -5.22694866595022, 
    -10.3697775665893, -10.8661435405664, -6.05533748614967, 
    -0.115990844370414, 4.42512947639905, 7.0617318768179, 5.57720718158874, 
    -1.22856703401718, -7.25133660196821, -4.38890777468485,
  5.324186773334, 10.7638084647545, 5.28523666180069, 4.48257892274958, 
    10.4117899099483, 7.59601726231476, -1.11628506805034, -4.92015012179954, 
    -5.87595470999816, -5.18324122114509, -5.53797199808407, 
    -13.3902947415915, -14.506257377188, 3.83248335490187, 17.5984269777707, 
    12.6406924680306, 2.07031653989326, -8.20890421591409, -13.6024703188098, 
    -9.34139044935997, -7.38952736662161, -4.54057080498675, 
    0.646254789483809, 1.43193142305978, 5.45887707543789, 13.1900036757778, 
    11.0223966135497, 7.96718492178897, 7.96378648070097, -1.01823679069239, 
    -8.35819428806321, -5.49907498387462, -0.384404034628509, 
    0.878486728677772, 4.56614910111472, 6.58760735847816, -2.29210012361724, 
    -12.1902363292883, -10.9101627731115, -3.43035718423223, 
    0.00562155588985162, 1.39405667853418, 6.62232732274148, 
    9.63189423898372, 6.0569531935516, 0.144270477824235, -2.32503898489649, 
    2.15145614587767, 3.36461206251645, -5.90493281227897, -13.1444288348543, 
    -13.0162110739888, -6.77711756195828, 1.91321285644953, 5.87769655252716, 
    7.16906844233398, 1.94483714695275, -3.33385355708656, -3.61151080142721, 
    -2.45062353303337,
  1.1975549874715, 7.03818654806387, 5.53933134303462, 4.43244007254614, 
    4.82475351749119, 3.82700239243794, -0.927406256031702, 
    -0.894770587286426, -0.764304317951982, -0.0935400448532807, 
    -1.47471420861403, -10.1714338645229, -14.8873297597856, 
    -7.33439670646672, 21.6759781913648, 9.32820674987845, -1.26755098042167, 
    -10.996211712289, -10.1264352564533, -4.76487759814467, 
    -8.44716913062961, -4.99232305472921, -0.0947791753732501, 
    -0.899914322121225, 3.28505416956978, 10.2702434285289, 13.07399235408, 
    13.612022449424, 4.60248094247989, -12.7312491911633, -16.4588649005268, 
    -13.8209436993621, 2.8374872198876, 7.72970664490702, 8.47750327916674, 
    10.5725332032756, 2.0055727243508, -8.35639840115466, -8.68199293615893, 
    -4.57396570256158, 1.32660231349005, 4.48329750911692, 7.06870600976459, 
    5.22103725416633, -0.31833646000283, -3.10017393696364, 
    -3.24816474992731, 0.32818229847182, 1.68355002871095, 
    -0.160384093997434, -3.72537527024945, -9.44401391089317, 
    -9.95219308678372, 7.23245586564813, 10.6626613619256, 6.66975234795836, 
    -1.32020756964839, -3.89460095915973, -4.47632512782093, -2.98822204877438,
  -3.83237234672392, -0.242234971521356, 3.99024327812962, 3.58650295850969, 
    -0.345044665464852, 1.1475705086675, 0.669293466262941, 
    0.178271744897631, 1.95498287121888, 1.14244972078849, -1.58609050982527, 
    -4.89383713819384, -2.09906179583069, -10.5611284127189, 
    2.63317335179006, 10.8193273395591, 6.55858055102598, -3.15562446431465, 
    -3.18803639411463, -3.34953809475501, -10.2308648721408, 
    -8.88269490909487, -1.18361685507944, 1.00672616966427, 3.33565854041763, 
    6.43275707122829, 8.80894003224421, 9.26265644953897, -0.708974354383093, 
    -7.39875290108771, -8.90576588261363, -11.6680386746181, 
    0.558843415111355, 8.40609008038024, 4.90066997903429, 3.79280411193326, 
    1.09868631000851, -1.40572383288154, -2.1923668671861, -4.52052528057929, 
    -2.64240474479519, 1.20414058340344, 3.72960648517372, 2.72438117037187, 
    0.157985557264551, -0.694003492288859, -2.0150476431477, 
    -3.92979117797533, -5.42520854322911, 1.97944689809989, 6.45446283709456, 
    -0.392824018298531, -7.15307230020351, -1.99722492039597, 
    11.0693039243126, 9.22187737695342, 5.17716581027575, -1.3787417035849, 
    -6.01150653928827, -5.44462294644965,
  -9.94724369297779, -4.37996251062805, 3.41101232048108, 6.78494792429863, 
    0.430521570798988, -0.364277927176875, -1.42246772176718, 
    -2.33163469690911, 1.65505653613015, 3.12091100951792, -3.29784954505314, 
    -3.500956103781, 3.75421258090882, 4.44971672908174, -5.68249200197557, 
    -5.83145747988155, 12.7523504183027, 10.9478973383845, 3.00815101012524, 
    -0.979424655882963, -6.75010012877929, -14.7640794059109, 
    -6.69294592841973, 1.24061169528306, 6.01929958447551, 6.83052973620639, 
    2.48928340445594, -1.68412182914558, -4.21626683527485, 
    -2.89004941734331, 2.09287378192728, 1.3741102063935, 1.55012525971997, 
    0.54205750003068, -3.42179237084594, -5.6144635131501, -4.99730288678459, 
    1.96983570702011, 4.97730976935064, 1.56075326287793, -1.8956749534137, 
    -3.39371860690337, -0.4064449824298, 3.25354947157886, 4.09760014750641, 
    4.451460915126, -0.363615789253723, -4.68417219375275, -8.89030887222866, 
    -8.97719381179614, 4.62630930560463, 6.39842566612294, 1.82800231401858, 
    -4.89580685664419, -4.43352246154103, 4.01687436681489, 10.9266474155208, 
    4.59463644955948, 2.26636219093625, -5.8323812190005,
  -12.1007409008064, -8.07710279986631, 3.38568451597718, 15.9221223689167, 
    0.0106459769305861, -3.66899019341629, 0.0680555136096297, 
    -8.42721360127858, 1.55574006306343, 6.46116786484117, -6.58913338651101, 
    -1.32771189047429, 3.58860766636905, 7.08441212030443, 3.7544197341656, 
    -12.2573243944829, 7.03068189667196, 12.3223924987773, 8.34298668755875, 
    3.02663860214945, -6.82485765314293, -12.3102748457069, 
    -5.19534351494817, 1.91259567704396, 9.3308582202006, 13.8199969285489, 
    -0.793737637546121, -15.6930697506, -11.3805770941719, -4.97610320469237, 
    5.00702428042359, 14.563127170473, 8.42334438165688, -3.59915172150987, 
    -7.05456554771927, -6.98094670132158, -7.24441708171573, 
    -1.01214277023952, 7.4267115561683, 8.58140243207939, 1.56413115928702, 
    -5.68360872278073, -6.95849898961285, 1.77049144521044, 9.57238574638882, 
    7.42760172432767, -3.95083458478341, -6.31726481792189, 
    -3.72295611847341, -8.34906455024241, -0.55455960569231, 9.4023748984359, 
    5.08510988561531, -5.41003967445815, -12.0440760449351, 
    -7.26932836494657, 10.2876534609014, 13.3158214754639, 5.94201556948032, 
    -6.24030248953981,
  -11.0167682732107, -10.965260086755, 6.39338281326439, 21.0541446593682, 
    -1.23738337896802, -6.35012614302901, -4.33173138528741, 
    -4.2930944481573, 2.74283166173994, 3.32386535763435, -2.67664083922628, 
    -2.16290098467049, 4.89253234956403, 0.17268427748832, 
    -0.165657742983827, 2.68836899614078, -1.93899198530153, 
    10.9883980572937, 10.1275789427423, -4.52803422659147, -13.39587398699, 
    -7.82986819379362, 4.15392146198349, 6.82229630411659, 17.6675140245769, 
    16.401214170515, -8.54469840593201, -24.422975263674, -18.0905085447014, 
    -2.4726123506931, 9.16562073483952, 17.4503884776271, 10.4029581416936, 
    -0.130104271990366, -9.24110235978809, -9.81224854926748, 
    -3.85379707852114, 2.02880593415247, 13.5670101451613, 7.06445889827203, 
    -4.61263080616295, -8.81185823712018, -10.0764794823827, 
    2.57084237202676, 14.8243103578399, 8.03687270117727, -5.32240685230092, 
    -5.58380634192843, -2.71567599604461, -4.00003664132275, 
    0.637553049206869, 14.6424021997828, 3.4754193775256, -14.2639374593964, 
    -11.7119588242618, -7.45327915022384, 8.43568349813647, 22.6699062321155, 
    4.23813430361593, -11.7409088230807,
  -12.3077442566777, -8.12067118093336, 14.1281724306579, 14.2338661463265, 
    -0.285719152407135, -4.8210849841411, -10.3463945603589, 
    -0.123865990016566, 5.33033376539745, 4.39163370744641, 
    -2.56382278741698, -4.54204573415382, -4.14134805783474, 
    -5.81607588762767, 9.32573326577854, 5.46772996157634, 2.90714259671991, 
    15.6897589780738, 0.9799966066648, -15.5422401384025, -29.5837480339045, 
    -10.7501178247187, 17.4045015685475, 19.1684344089282, 26.978909132044, 
    2.93266965542676, -20.4099903683219, -22.3944060855082, 
    -15.0412034162306, -4.41250996166811, 12.6002208849748, 21.7832818430293, 
    12.3541361565616, -5.27148085758242, -9.47838225992006, 
    -8.07907273144419, -7.47613728037161, 9.95076859733875, 20.4770684560086, 
    3.7876473192902, -10.4599791898725, -13.8566049394947, -9.7931898855234, 
    7.48086729285762, 18.8322649435984, 3.48418141514862, -8.06670995003124, 
    -1.08518212219702, -6.09692879588981, -7.77539196890365, 
    11.8613931285035, 17.1943497448248, -3.32029670156769, -15.8059045844449, 
    -16.203222605015, 0.279905353966314, 17.1039643611174, 24.5442322715411, 
    -2.99957747407745, -16.1755533153509,
  -8.79767720627783, 0.218565952167803, 13.7037357592568, 6.3736294256032, 
    0.524966047987127, -0.282422192914917, -9.54134440267241, 
    -1.15331734513919, 6.83098617706792, 3.22574239206665, -10.4273103879117, 
    -3.59895883096013, -7.3700982980933, -4.54303046628811, 11.4947948577383, 
    8.43668616097893, 16.4493253074536, -0.996121003551056, 
    -18.7569348478768, -15.2794164583393, -18.0697738595681, 
    -8.84452342904632, 16.1808546642856, 30.0178318493135, 17.1031732921707, 
    -14.6478336397791, -21.8367902127853, -16.9787717250089, 
    -3.77763819893912, -0.00662141400348904, 13.3835349829975, 
    13.6269394027077, -0.642356254409575, -8.40243196163041, -4.193507989787, 
    -4.30808610677338, -4.30088926803516, 12.7683076297139, 16.5271786312508, 
    2.61335476132677, -15.682167261567, -10.8855592276546, 
    -0.154445809253625, 11.3329901877916, 5.71449968810403, 
    -7.37352543214837, -6.75342270165781, 1.43789697128802, 
    -5.95460363062229, -4.68060797119433, 16.4242997357379, 9.65181392124056, 
    -11.3866856503007, -12.844183234952, -9.1710383650629, 6.23655982255927, 
    19.9427994929346, 9.40876500099497, -8.91032504819749, -13.4484958765226,
  -0.310660429476216, 5.35305218485697, 10.461356905953, -3.35713075589296, 
    0.399814241941464, 2.25381108616324, -10.2993798193308, 1.2743879183676, 
    12.0845593165163, 3.5420746586551, -11.7200982759968, -4.12721240224286, 
    -5.04056558774798, -1.5705637116855, 5.8687924641041, 11.5002586255022, 
    -0.779795489793761, -7.87890693006295, -13.9567351833658, 
    -6.30238521441671, -8.61057560323691, -0.124004977182193, 
    18.3095139280114, 21.5804162680536, -0.49767876819771, -10.9654674130933, 
    -10.0514895477584, -1.97857968263305, 5.7433508221804, 2.90731381335532, 
    6.01454462725263, 2.00008365518113, -7.22525070238379, -1.46889134632749, 
    1.63458203873611, -1.52585110080124, -1.20673650465024, 1.76473164991414, 
    3.29452610688251, 1.17171251033247, -3.61592852801724, 
    -0.198315307356127, 4.57233180145733, 1.58956816471683, 
    -5.12254384837831, -9.32854011921062, -2.40820172514733, 
    0.811138437784209, -1.12736326972008, 2.2297343607607, 8.65738098172328, 
    0.433718663511723, -9.37472949256382, -6.00610315588907, 
    -2.51705917414357, 5.51542868952105, 8.18795754243468, -6.96162382750676, 
    -10.2593120693593, -7.64078453695672,
  -1.43618973280492, 4.89080130512867, 7.63728951602956, -0.878891411920541, 
    -6.55660651611578, 11.4171509391861, -5.47795569897624, 8.02150030018387, 
    25.9514708709356, 5.1661791385163, -3.79466973368118, -2.96275577331359, 
    -2.25231281144494, 2.4115129554706, 4.64090886462556, 4.9535795650645, 
    -4.02099372344019, -3.38055869674623, 3.68905268513334, 
    -4.37709184870448, -9.04893230051642, 0.908646224694664, 
    14.0243428285207, 1.97440348050911, -3.11556815128194, -2.71491259134984, 
    -3.79407082220187, 5.24925134483026, 1.24935805485798, -2.06921880621403, 
    0.644619095984029, 0.532080135402306, -1.82702229801675, 
    -1.56980349815275, 0.75194101312745, 1.51405433707447, -3.07160299913523, 
    -0.224140004046534, -5.23798586670094, 4.08948052877195, 
    12.6970527642344, 6.851939637472, -0.937470328512956, -3.97070310663839, 
    -0.38995631559597, -0.222077439873251, -3.51925230743456, 
    -2.72799439379883, -0.176306814047797, 2.103444096987, 3.37835248695372, 
    1.48151912569824, 0.541287102014514, -1.50230230858049, 1.02409883192597, 
    5.73870667595568, 0.245820890337054, -7.74342969080525, 
    -4.24063595014993, -2.52891415312776,
  -2.33651982923945, 2.48192970827806, 6.88083025693474, 8.17470975925422, 
    6.27785013250933, 13.2537240561707, -9.07626283396818, 13.5666878001114, 
    18.5801514290991, -7.17826400375516, -2.16849928350376, 2.57808734195953, 
    4.70032312415608, 5.89204580762529, 5.47400934020017, 1.57044757173872, 
    3.06129240715795, -5.1441489805563, 0.781377926839922, -3.26532104378459, 
    2.24521444756595, 4.86323968349095, 7.18184175170303, -5.99521998200766, 
    -5.78244873873405, 3.41237824066236, -0.801499852171684, 
    -2.71163187330357, -4.16221842176187, -7.10372740289578, 
    -4.17352302848491, -1.62035099585428, -1.29519750294514, 
    -4.40629009927743, -3.11040965430857, 1.26429409377626, 4.52036417231322, 
    2.22779203764313, -0.820374349489864, 2.33257383165089, 3.54448363728581, 
    2.32733314488818, -2.08609010977871, -3.43864725218456, 
    -1.83298455090056, -1.02324326457193, 0.97446749210995, 
    -0.166750707739925, 0.212441970904651, 6.50977024621715, 
    -1.75630970151681, -0.721811783928522, -0.917620382074002, 
    2.65605923549823, 1.17070157222872, 6.1126411388487, 0.155652527394471, 
    -4.97514916941484, 1.6901168730788, -3.10752407071206,
  6.780583154506, 7.16368452201328, 2.52878689663383, 4.26505337098219, 
    -0.685156648197058, 2.04442620445053, -9.93452205428011, 
    -3.78387637032764, 8.59116107159305, 3.54180394981366, 1.47259429935605, 
    -3.97055701464355, 0.89142537334879, 6.75248114176602, 2.08945849231013, 
    0.907705260127619, 0.526759528259366, -1.16727863505379, 
    5.62399668987231, -0.243632341430088, -3.83996860123064, 
    2.27971649009146, -1.2406920885697, 4.76375359283847, -7.78254219412533, 
    -0.866744683888403, 5.04587156050388, 3.59882778925228, 
    0.305309293345339, -0.329603064482657, -1.63467836965215, 
    -6.75057292975724, -2.01590652441221, -1.6003477905227, 
    -5.05785767413807, -4.6055142935725, 0.215285447357467, 4.49489636041416, 
    2.72652612426963, 2.45638588745295, 2.74636428838812, 0.421808210516128, 
    -3.98657006689974, 2.32372525635535, 0.96578710416494, 
    -0.242984081267983, 2.39347413759487, 3.74097624158473, 2.90534948640887, 
    4.59158051729818, -0.663947343685256, -1.89780145918883, 
    -1.70595659176174, 2.78896728309596, 3.00952726603319, 0.785627627911235, 
    0.503952381692132, -1.62044377561413, 5.75795446762405, -11.2665851013789,
  -3.43438901082069, -2.46923895152038, 2.9554251744205, -3.33571556889156, 
    1.52088932603299, 4.056074656381, -0.40761842841463, -3.49076762349046, 
    -0.369284599118763, -0.269496368482037, 6.56840658711229, 
    -0.287806794390103, -6.68781582879313, 2.34137810001309, 
    5.77800450271564, 1.1248232617842, -1.03134999676785, -2.87698315281094, 
    1.57982751987572, 3.49968865638464, 0.632936928764725, -7.46167740585724, 
    -1.83949667633621, 6.69938489239569, 0.523434493878388, 
    0.387624490291425, -0.36184588735229, 2.46132369854509, 4.26889216210873, 
    -5.7539370638274, -11.4344144273818, -0.000310767306037821, 
    4.10435291515578, 0.293646965921842, -1.05108167365512, 
    0.587603721042563, -1.51446056447336, -2.81785659280632, 
    -0.006026686471425, 2.22142921697594, 3.52086944677762, 3.09471110085431, 
    2.40303386103197, 3.75388367529904, -2.6729677375196, -6.09613865810488, 
    -0.389620002055043, 3.38840296838241, 3.72820716721841, 1.34519025601807, 
    -3.00961318833376, -1.57490405749068, -1.00826009227856, 
    0.732996676008638, 1.86107369482263, 2.78805098294466, 0.830580815787736, 
    -5.07196955080392, 16.2908402955412, -23.6555783212225,
  6.80155065622094, -5.96379310077859, -4.20300785046729, 0.139364650519265, 
    1.40038082262412, 4.31384941898723, 1.87667469765658, -7.58372482428907, 
    -12.8726214004978, -3.44482547752895, 11.683125647768, 10.1033282142348, 
    -7.97047154894853, -5.34678388024887, 4.28075560617066, 5.29155539874912, 
    4.17171251565099, -3.10873590246774, -6.24596488575965, 3.3334905717335, 
    6.90281772586279, -2.84445975970761, -9.03185691663438, 2.64175978831936, 
    4.35178264927132, 4.89506370596721, 1.19764549859987, -2.82450396855642, 
    0.151351326086094, -2.60581018228139, -10.2716531258339, 
    -3.76967511397524, 14.116108780173, 14.714480073979, 2.49632711842815, 
    1.21665795121243, -3.89788419369461, -14.0428689607478, 
    -12.2781732474696, -2.78852030520789, 7.56751081488565, 10.6243024939315, 
    6.45483797413457, 2.73284578708801, -2.00046479224852, -7.29731261484431, 
    -7.62360880903824, 4.91981843079038, 8.59286739845475, 0.578744078842846, 
    1.74233537192996, 4.54922179044244, 0.0201807299638734, 
    -0.0951847466472608, 0.632978087750016, -1.12877662020518, 
    -7.37325017672913, -6.21837978348202, 16.982001620906, 0.157249925161029,
  12.8231004344166, -2.90746705524184, -13.5646107131382, 4.71191464036963, 
    7.56442572171103, 5.40108684280472, 4.71903547699375, -9.31438878702908, 
    -25.2305358263736, -13.3465146509209, 13.4557898772631, 19.8934346760864, 
    2.09287077926268, -5.72530870591185, -5.01095191807839, 
    -1.36832622332921, 3.90829149250398, 2.38456440439671, -6.46151800328032, 
    4.33956673909414, 6.91409414751413, -4.41225155593883, -9.97364542377507, 
    3.51785947628569, 8.1807326817756, -1.32939216867922, 0.75933992208076, 
    -4.08758326236439, -3.44281324237689, -5.03425778664329, 
    -2.33438677608747, -10.8357065000384, 9.12449660027986, 24.4728913348774, 
    13.9987843138188, 7.48905829698459, -5.04637292622819, -20.2981409976658, 
    -22.0181923366578, -11.1494727712119, 9.37778565144819, 16.7530033657245, 
    11.1451577132538, 2.01274515867951, -3.71302663101005, -3.24149552716281, 
    -12.8614426601128, -4.94406815019329, 9.30289698336932, 3.84305269272728, 
    2.69184116062484, 10.0739221496531, 6.81033952195613, 1.26563783314163, 
    0.151139084079854, -12.0558651465124, -17.9866291091972, 
    -10.364623081681, 13.9330803440029, 10.2371484710617,
  6.65377126435651, 0.698569879303124, -10.6262259850054, 1.88855945684777, 
    13.3665047992521, 14.1219067400907, 7.20524352885079, -10.2466946983817, 
    -25.7345855955061, -23.3621038148689, 6.03955484008842, 21.0474294213717, 
    14.2182919965212, 5.67834657168551, -8.69164214644203, -16.7545497588563, 
    -6.90155404714178, 6.56133137861561, 5.33883192690022, 7.27743745744496, 
    4.80624034923832, -8.55066733617567, -14.0875900085923, 3.33119968946237, 
    14.4195622835784, -4.08272912348909, -3.71329344170217, 
    -3.62315575605834, -1.70156939884536, -1.13162452076467, 
    -2.37408960953549, -9.77726920836335, -3.37343459097995, 
    18.3917050194229, 21.2802757540283, 9.10910489100316, -0.76301555323053, 
    -16.1201380890134, -20.9611205320022, -11.9061462742401, 
    4.53811275876416, 12.0825564262773, 13.3200793878155, 6.38613153376059, 
    -1.4422935028935, -3.02376424972528, -10.3051067214448, 
    -12.9901333886966, 3.8926641074925, 7.23499281334582, -2.1498253918901, 
    5.56891540641575, 10.4608861545018, 2.82063668720387, 0.280862662491332, 
    -11.5255373190383, -15.9002309539248, -14.8001075580392, 
    5.81752206379209, 15.5756284880613,
  4.43308502464666, 0.603715056483948, -4.79249518306659, -1.91109645890112, 
    12.5943940795462, 14.8453596746268, 5.69520835348362, -9.30686525752282, 
    -16.9701791984699, -19.188911012007, 0.904914890700067, 20.992679356458, 
    16.6383712618477, 10.626551810535, -6.73589362413514, -20.3209550172758, 
    -13.2847149518492, 4.27228899744155, 11.9791485685508, 5.78708342445745, 
    8.16085198271909, -7.4069139087579, -19.954387566493, -2.97400247699097, 
    6.73033287198882, 7.88471412984914, 1.22545623386585, -5.19373218378611, 
    -0.441187339200285, -0.842207227037084, -4.43852243017759, 
    -7.90988249411874, -7.80123146684565, 8.68438325441277, 15.9875476885745, 
    11.008450031865, 5.98639006031044, -11.9069262147933, -18.5462988348972, 
    -8.74314043444384, 0.836024276333134, 6.45238182394427, 11.1939967411704, 
    8.37244215208438, 4.72531470082901, -7.29741600680734, -7.96367483060413, 
    -6.62056889447806, -1.76696287464561, 0.378163956943193, 
    0.28248790350049, -1.30349722997124, 8.10734961329688, 7.15461245042262, 
    -3.29778216747723, -3.46165809867532, -8.24128495781176, 
    -8.43429024487935, 0.720993814537463, 8.60180022146396,
  -1.51720678937265, 2.63386023294224, -2.4304549476621, -2.8557480488586, 
    7.81562521611004, 11.5637773692638, 8.97906845101186, -5.14728751929709, 
    -13.0703613195212, -9.72019234159042, 2.48320088342379, 16.420951707814, 
    12.1841790677162, 6.02614707363284, -4.49706501604936, -12.7901293694263, 
    -10.154157409643, 0.174861878477531, 5.61918481764732, 8.01828738211493, 
    7.1953360189408, -10.0140762588168, -14.7197099111075, -5.21283330439456, 
    6.11849172681273, 15.5343747913608, 2.7369646216761, -0.894669927667079, 
    -1.528322836298, -5.97000250234613, -6.98199837021109, -4.95734725759443, 
    -4.54690485631127, 4.57408140768106, 12.0155367439943, 13.5621373444767, 
    3.31747606602915, -11.4336959937606, -10.5703631794261, 
    -3.02338096446373, 0.814235067086741, 1.56230226915702, 7.21350018118118, 
    10.8767600042805, 5.44943751537318, -6.78874270556847, -10.5700451762087, 
    -7.60077084787981, -6.55190188921204, -4.68550966693615, 
    -0.0561615402943071, -2.54827396708002, 5.31212544910804, 
    9.57800062614114, 5.73439255189137, 7.9140724123552, 0.131742684593951, 
    -10.1373544787306, -5.90209492487801, -6.23333363019205,
  1.67482452531817, 4.10471759653408, -0.967831007386572, -0.445460742484134, 
    5.78294823322613, 8.48042618743781, -0.814535729141265, 
    -7.70020876129814, -3.68313886574883, 0.590196290386365, 5.7732404483191, 
    8.55033404274664, 5.67623305311711, -0.530432169463643, 
    -3.18793464600043, -6.8674971214044, -6.44405805962551, 
    -0.876698617551269, 1.83936242395845, 2.37429531837793, 
    -4.79753791940808, -2.00571475110371, -0.204295166398505, 
    -1.74318558209815, 10.4448327768814, 9.11336783263432, 2.46345480236423, 
    2.70889438573005, -5.62982619222488, -3.37989087031622, 
    -3.66139892485428, -2.90223922296091, -0.498705670825593, 
    4.16451595002799, 6.07460958989183, 2.81363692188521, -5.45957418301792, 
    -8.97068156044517, -1.10997452680729, 2.84780158003298, 1.63498849436664, 
    2.10406534689762, 7.45113917349209, 9.78336844053275, -0.897747740715898, 
    -7.3452800109551, -11.9703102139225, -5.60673592872626, 
    -1.68805196022532, -5.47896307846065, -0.54189125066885, 
    -1.85211161891162, 2.94667253770138, 11.2421978152504, 14.5203732301268, 
    9.05631553116211, -1.30561065436697, -10.2970208422322, 
    -8.91734681859819, -7.42519292132275,
  10.5600993165872, 4.37172078536821, -3.1122123619055, -0.983782951185424, 
    2.12454508826395, -1.75444550181655, -8.59492632731437, 
    -1.88237739389817, 5.30775416207339, 4.3629747005995, 4.39249097327283, 
    3.47975852149025, -0.43240135718596, -4.17946956323919, 
    -6.38396662618075, -9.49716908260007, -6.57703538563703, 
    0.956910320116374, 5.66809821862262, -1.32408127051535, -5.2704373811578, 
    8.55933548335627, 9.41957907006124, 1.58407355372833, 2.99076079901859, 
    0.938460977030132, 2.0483669188028, -0.819965348488466, 
    -3.83711657824524, 1.10407064644535, 2.2460796162618, 3.46490319085207, 
    3.27231665615141, -1.87561129659647, -3.82834582863339, 
    -6.96439277810975, -11.2070867551898, -7.83020895090786, 
    2.56352838220803, 7.95765527769155, 6.11995407246015, 9.37508467469205, 
    8.06760721346736, -0.2941150596348, -5.86203066229322, -4.3012641211098, 
    -3.74638829250691, 4.85729249005391, 3.62195615423024, -12.2585001175877, 
    -4.14491765060896, 0.908114983404523, 2.69079743600393, 4.63094883084592, 
    3.96450530060492, 4.70155413725368, 2.16801954497412, -4.7815134845602, 
    -8.12209699221533, -2.0899217885519,
  11.1280390247505, 6.81046939933924, -1.58399515503101, -1.00990295476897, 
    -1.19278897305734, -6.06747351889798, -6.97875729348458, 
    -1.43398111164835, 6.03703593413785, 7.35994262088482, 3.8213196198282, 
    0.581791488543972, -2.49878080090241, -6.02322404734054, 
    -8.85003831893953, -10.1547510435658, -6.8654886918572, 1.83045002053511, 
    7.25376875372804, 6.42777755687422, 6.76815427604056, 7.03218041885315, 
    3.12609844792499, 0.593874672272016, 0.573303911305631, 
    -0.157458158381473, -2.51715744612844, -4.85818001249952, 
    -3.34032859985961, -0.0857942669918578, 2.9465965735754, 
    5.99612344823283, 2.62780327853782, -3.32693967658662, -3.70466076734948, 
    -7.03986052852216, -11.8626379482384, -6.85937350361317, 
    5.03243628365108, 14.7910239241784, 15.7811770556726, 12.3963706330412, 
    4.80040711757204, -4.1202128650548, -7.27695762681857, -6.14376166952724, 
    -0.391604072006802, 6.65905187715975, 2.5750942033417, -9.05007239853831, 
    -8.97655422889551, -3.52561073526222, -2.71363836850319, 
    -1.62429899609222, 0.356830059360316, 2.35752864880493, 2.28382637947481, 
    -1.73083378912275, -3.93935002582694, 2.5225472825103,
  8.86829578489544, 7.30842679467364, 4.47025553672674, 2.01336213349285, 
    -2.05167397737459, -7.95174151659696, -10.0730359348937, 
    -4.68349797189595, 3.25303658754586, 6.95766497946276, 5.99575857380624, 
    3.66443058034665, 0.953601094220854, -2.94643081420099, 
    -6.84901253842493, -7.59200344059472, -3.91211017535616, 
    2.20777998188836, 7.06889267437151, 8.21211060662937, 6.50315662500961, 
    4.44402555335636, 3.69680493149982, 3.91012479499768, 2.96562684393616, 
    -0.961185573910527, -6.55370652231898, -10.0588020846246, 
    -9.23972615828524, -5.53338211182898, -2.48477730946825, 
    -1.58269194114628, -0.583493863736683, 2.03222465473443, 
    2.46752764025258, -2.18475422348837, -5.64766347875491, 
    -1.08845461275788, 8.32141815361648, 15.9921127867211, 18.57850370022, 
    15.2349521256353, 7.69205669691247, -0.673870962405759, -7.7885122897192, 
    -11.8839082383279, -10.1995133367923, -3.35019579044502, 
    1.70872121231577, -0.763698556193874, -7.3581737450675, 
    -9.38341950615108, -5.30713254304977, -0.944918276179371, 
    -0.158774217251893, -2.1113631374418, -3.907452952029, -3.00901406806686, 
    1.32600730215763, 6.5354977945707,
  5.09654024286252, 6.76571534221355, 6.33527659159213, 3.9970797131073, 
    0.0580590273221122, -4.35860535372469, -7.29449536269939, 
    -7.07791426150549, -3.63551305313294, 1.14191601636649, 4.81087603988048, 
    5.77124784962348, 3.79848404808811, 0.32517092589755, -1.99724303313544, 
    -1.12954412030845, 2.49691658040757, 6.3278330802254, 8.16612231761206, 
    7.75775419124389, 6.49995629832648, 5.92753257881556, 6.22675133313313, 
    5.90053438190979, 3.15076529539984, -2.19458980062951, -8.24944767082484, 
    -12.5326952299979, -13.7757852218563, -12.3296140646687, 
    -9.18566437288555, -4.92846593741496, -0.0549402716413629, 
    3.90757463901111, 4.91490519267706, 2.82789851317227, 0.264957492175581, 
    0.488236815331767, 4.28548094168898, 8.96199283071482, 11.3550872772558, 
    10.2889412601869, 6.38492859472461, 1.05763846057601, -4.03308726121271, 
    -7.28212411566082, -7.8281865251891, -6.02004827097048, 
    -3.26391557662643, -1.27361017793914, -0.61007638241195, 
    -0.541294291396608, -0.297599566776526, -0.454742158073858, 
    -2.19806773947897, -5.24979592122852, -7.53741401801721, 
    -7.00410333915823, -3.45486635533018, 1.32958981386604,
  -1.70964914333507, 1.11210578701888, 2.9360686431048, 3.20175246517757, 
    1.99850759012491, -0.043264761830017, -2.02591172445034, 
    -3.15928593343619, -3.05538939280394, -1.85437356473009, 
    -0.224761915809722, 1.06509067455361, 1.68024243219764, 1.87203556520016, 
    2.2139038701715, 3.17939537521034, 4.8002664906399, 6.5911318914519, 
    7.86111065191457, 8.19168788460797, 7.56517819831457, 6.22774963744783, 
    4.42499262479391, 2.24528926735857, -0.329469607414148, 
    -3.27282596564171, -6.33257406199719, -8.94849937656891, 
    -10.4191830132177, -10.1684419888346, -8.00450395354532, 
    -4.39357260791098, -0.411627301347247, 2.71365438840399, 
    4.16335490706996, 3.85329310009105, 2.42682236607998, 0.822570902627761, 
    -0.18147241190457, -0.19812678509726, 0.522379091886742, 
    1.22803443080737, 1.25882246854643, 0.471780627913666, 
    -0.719043202494768, -1.66368553120875, -1.88297545973968, 
    -1.28308579984018, -0.0625165679828535, 1.39213840904991, 
    2.67972919651385, 3.45623635827985, 3.31338403440387, 2.03658143843346, 
    -0.182674805356393, -2.81436276674956, -5.16290154220284, 
    -6.51405243762438, -6.32386438430584, -4.52863782317413,
  -0.830942909007372, -0.68977260871087, -0.468771252369503, 
    -0.216644510564877, 0.0200104048380254, 0.222044142301965, 
    0.375135391929922, 0.467785566995632, 0.502485853892534, 
    0.494549951490028, 0.493148304569599, 0.551870545149785, 
    0.695991218810392, 0.918574319871883, 1.19497317915357, 1.48516278689069, 
    1.74466256232481, 1.93785248110497, 2.02574290778099, 1.96080480408685, 
    1.70911094650212, 1.25556460635859, 0.623006570070456, 
    -0.132664620932614, -0.93222554918056, -1.67368742771848, 
    -2.2644567828659, -2.63771999571281, -2.74368386604998, -2.5701937594754, 
    -2.16903216087145, -1.62150541583233, -1.00783874462876, 
    -0.409584823524948, 0.0902507486505314, 0.434719136372979, 
    0.597072954328891, 0.581695071820981, 0.431001186337763, 
    0.207649130538047, -0.0223699268647248, -0.18611249452731, 
    -0.230216030003615, -0.148247901846373, 0.0211004414973903, 
    0.224830630597154, 0.419614819233677, 0.578120594031707, 
    0.681148737274401, 0.72546651443892, 0.701678489758768, 
    0.580854366412161, 0.385280445238711, 0.151368934619055, 
    -0.099372820953807, -0.330049004488905, -0.516386878228678, 
    -0.674196093395887, -0.8031679010168, -0.866194039755007,
  -0.920165223119996, -1.9606260229677, -2.94249723453981, -3.80143530871806, 
    -4.46525690046493, -4.85624930322331, -4.95488917655344, 
    -4.8026962805427, -4.43692736678313, -3.90023662712362, 
    -3.24392129840348, -2.52630804669138, -1.80168414473207, 
    -1.12299992145145, -0.526159860659726, -0.0203936273938838, 
    0.390029850055706, 0.68250095381592, 0.862053430921432, 0.97113698490228, 
    1.05459521341048, 1.12603940350096, 1.17743994038336, 1.22586610577757, 
    1.2966599167856, 1.41881924586872, 1.60906948949856, 1.84276068425561, 
    2.04144560360104, 2.17354493372664, 2.22976246109388, 2.15239563378512, 
    1.91928975407908, 1.56199240783269, 1.10933876374311, 0.583787167093737, 
    0.0112635858907869, -0.570566646327162, -1.12191649708666, 
    -1.59787845525327, -1.92949156527854, -2.0690411487718, 
    -2.01112649873649, -1.76801609877246, -1.35194820883616, 
    -0.775878613175074, -0.0603782216283259, 0.750284556398804, 
    1.59031152950089, 2.38050494801121, 3.05625106268128, 3.56345231478893, 
    3.86276185912513, 3.93664207904511, 3.7740588000315, 3.38981666786076, 
    2.80687327770223, 2.04980750410451, 1.14579961263143, 0.13369088793373,
  -3.61045074510779, -4.06460969039647, -3.67406120635378, -2.68609030962766, 
    -1.60367377761822, -0.936071309598789, -0.844710444126519, 
    -1.13740785910817, -1.61622969335897, -2.14704307475856, 
    -2.57427886535092, -2.73746429593239, -2.55461211963148, 
    -2.0134561102584, -1.21316397397343, -0.3595981697364, 0.326111473798985, 
    0.770467234499443, 0.882250045734146, 0.68938246477603, 
    0.477240980617616, 0.581301648890354, 1.2122912975963, 2.28047095632303, 
    3.44298620492447, 4.22960054251047, 4.2971319968624, 3.6395477574796, 
    2.64229237091572, 1.71102870750128, 1.16185782849842, 1.26624855505712, 
    1.93520175872931, 2.69900751228364, 3.00730443293536, 2.45073219527723, 
    0.924548099029559, -1.33542796880953, -3.77990606822738, 
    -5.75471507194324, -6.79493538747346, -6.67507721701294, 
    -5.39323696434354, -3.21741696006833, -0.619459806058921, 
    1.90279601427583, 3.89173223442878, 5.00451821870536, 5.13266336445147, 
    4.44710119231961, 3.29569419753236, 2.10111682632793, 1.21180498355986, 
    0.807376639467948, 0.853851107558422, 1.02102977328001, 
    0.889237475621543, 0.185206041312071, -1.05155342592494, -2.46975293767415,
  -2.56703176783057, -0.473695924451997, 0.80473781852619, 0.828183056243411, 
    0.788050638108534, 1.83215037260683, 3.12929717099395, 2.75682879986318, 
    0.307043466352694, -2.74002494835475, -4.83859119024437, 
    -5.52175660323551, -4.93263852936798, -3.36461792946383, 
    -0.808878790397017, 2.27993312684093, 4.48249342835775, 4.30799520442401, 
    1.93517492497787, -0.526293769150145, -1.20982516052037, 
    -0.405746879058384, 0.565974497231589, 1.3927640042472, 2.65279098840831, 
    4.43150190151587, 5.58768984316832, 4.73062628173028, 1.54013135563607, 
    -2.12706581051834, -3.33265725891808, -1.07944089674969, 
    2.81170758253582, 5.49584828106263, 5.24869528623399, 2.44531453058149, 
    -1.18313245919276, -4.1883436874036, -6.23756554246972, 
    -7.56746908756346, -8.02184006026288, -7.09238637658178, 
    -4.52506750186967, -0.835953343027665, 2.66764830355795, 
    4.67492751284241, 4.80783375738243, 3.73645143368174, 2.37104441447039, 
    1.15318822747737, 0.240171790536341, -0.193394673804843, 
    -0.118795294688607, 0.305545708661468, 0.67862002286698, 
    0.649697295678742, -0.0696775310114948, -1.56500911041302, 
    -3.22404240220555, -3.79607720064604,
  1.49959723321405, 6.40781287050771, 3.87117117277931, 0.261028743166042, 
    2.40426253117112, 5.9948748099599, 5.02199081005069, 1.8611262809082, 
    -0.493034319917173, -4.11298139764482, -9.3233492280333, 
    -11.6342207456724, -9.27271714025076, -4.1416905842927, 3.02097436218076, 
    9.08162625276137, 8.8489832159387, 3.05538263118392, -3.15971730350394, 
    -6.01990314285204, -4.91176293498784, -1.77528118190116, 
    0.259374941092372, 0.702513730597368, 2.99348654376659, 6.88095107116368, 
    6.56816407649186, 1.0147980137194, -2.39491441718846, -0.703125206468271, 
    0.72701949134299, 0.0940940032379843, 0.730628328564417, 
    2.67998802002198, 2.6582829674773, 0.40912730732026, -1.74211283911466, 
    -3.5107378948623, -5.37562762780385, -6.40084850185577, 
    -6.38201109822329, -5.26394570631182, -1.70086334664751, 
    3.65420450307542, 6.57044980069918, 4.92982904897034, 2.17293900634186, 
    2.26827762860504, 3.57776022803209, 1.42457657724062, -4.3355755821152, 
    -7.66369150568242, -4.98650158170275, 0.34239815266426, 3.55728808740328, 
    3.73939098237236, 2.64799013434821, -0.462492123532356, 
    -5.08837321600083, -5.13540555841153,
  1.878041049097, 7.15911682377812, 3.28373342470258, 1.26344972059062, 
    5.8356826797258, 6.96889484043604, 5.95674432221081, 5.06449569554201, 
    2.26690210123229, -2.93454864873998, -9.48448317948973, 
    -14.1184060950716, -13.012629316849, -4.06491163944673, 7.75635896075959, 
    11.5029382565541, 6.23880101958541, -3.30469833304153, -8.29120386144359, 
    -8.11309931280021, -9.42251003720286, -7.5584847121883, 
    0.301790432865508, 2.88508981558766, 4.10127419272333, 8.76128531641773, 
    6.58478563469008, 0.751698047736165, 2.00228023452693, 2.11935514146138, 
    -2.27804772777895, -2.93039333150757, -1.00729842498029, 
    -1.06190488354878, -0.0876624672440554, 3.89820111664193, 
    2.89724939950262, -3.73562020853124, -6.19107720406915, 
    -4.48316606371409, -3.6091691627044, -1.49105624998344, 2.55913381261702, 
    5.7923638304584, 5.87327437216011, 2.6165543577439, -0.00386424657926438, 
    2.21508103801376, 5.63002913517477, 0.552530601991467, -9.52575681162718, 
    -11.4694833315793, -6.71326401990319, 0.0711145709480117, 
    6.04184941341579, 6.57079435882006, 0.990895852757069, -4.28644619828685, 
    -4.44406498280868, -3.25005411931892,
  -1.68199963049346, 4.6311388379529, 3.30397267064567, 3.44562248167856, 
    4.59543847978134, 3.15463728079666, 2.93305869031551, 6.69812105127305, 
    6.25658725249141, 1.45770107966588, -4.81393221727953, -11.8620883550363, 
    -12.0959462263072, -10.3946618523948, 12.1946913599108, 7.6028999409986, 
    2.24586204825026, -4.23848827228344, -2.68145638902207, 
    -5.93129685634677, -11.1386118263715, -12.0586658382729, 
    -1.72040924523533, -0.640487774953174, 4.11528172591051, 
    7.21722892703122, 7.090987865426, 7.72646744748913, 6.32995284734918, 
    -2.65317532098428, -9.97801100378405, -10.4802035104617, 
    -0.652931167362286, 2.75661865003613, 3.01902762200059, 8.62156907910722, 
    4.46948041976177, -4.32920366017541, -6.580002298631, -5.16002678901811, 
    -1.58489605758081, 1.60852655456268, 4.76789900227765, 4.66196720245422, 
    2.65481084988728, 0.230421815723215, -1.35083088637111, 
    -0.428841405543423, 2.32019500336902, 1.07889101792456, 
    -3.17570883173952, -8.20853880339608, -9.49137640469157, 
    4.62393130147853, 8.19976252899175, 8.39737559831418, 0.986903134342792, 
    -4.03118034068909, -6.35872607452224, -3.24285443898995,
  -3.46253869843325, -2.40513637592049, 1.27183220115739, 2.40063938224098, 
    1.03429235227118, 0.467672601246483, 1.20930177677768, 3.69650553097095, 
    6.18563872235044, 3.33074742370961, -0.727798578653113, 
    -9.41037143033752, -1.45928607452841, -8.92873961721129, 
    1.13330434462507, 6.72278952439121, 4.37653199990569, 2.87789157830924, 
    4.58178907973539, -4.0057482540426, -10.3790818009315, -14.5673746978548, 
    -6.40366290776128, -2.7009425959055, 2.7393574012179, 5.15313571616031, 
    7.87507315876414, 9.7429705219504, 3.8726581275736, -3.59596545003031, 
    -7.44573401421165, -8.77406308302161, -2.77670272936346, 
    4.64605391680111, 3.49563325105486, 4.62455879768969, 2.40622688801856, 
    -1.79288370854455, -1.47277609911379, -2.75440572682955, 
    -2.75000930911673, -0.418807185685646, 2.57141726866256, 
    3.52996194961762, 3.11058968034729, 1.51515881445607, -1.02946556230026, 
    -4.0835110693053, -4.27244846346532, 0.919584866503336, 4.48121327435951, 
    -0.122715288623321, -7.92181118704275, -2.95820093763852, 
    8.75814641767841, 8.18455948390882, 4.53170165522112, -0.635564821980641, 
    -3.7831469172354, -2.50599619231176,
  -6.66426767202049, -4.88720837870754, -0.747981393108052, 3.75900783662211, 
    2.40269386312068, 0.576452117413538, 0.0993756623224665, 
    -1.6410562547864, 2.11977477268603, 2.17298993985281, 0.868636941410923, 
    -6.20245796750413, 2.29066825589412, 4.87657272696449, -2.91090845047037, 
    -5.35019730899639, 7.03116143076869, 9.24651718702321, 6.84077970115501, 
    1.4151578263717, -4.71192294133309, -14.9059610482393, -9.74251099639604, 
    -3.1121785754335, 3.92872078045612, 5.20989742730022, 5.22588646133503, 
    3.42223125864713, -1.29769239418142, -3.09663423094897, 
    0.414476149496493, 1.39502333665956, 1.60912250061644, 
    -0.190284368031256, -2.33554372847368, -3.77686695661427, 
    -3.38444517479823, -0.681893040110225, 2.46670373689642, 
    2.37880032213416, -0.241323827725851, -2.25617298854816, 
    0.137810052183296, 3.49069251071473, 4.44783498518827, 4.69338687045547, 
    -0.0498156962241839, -4.36055493233503, -9.17478156971337, 
    -7.19335627716598, 3.5401970449611, 5.77192650347878, 2.89213217727909, 
    -3.20527876903975, -4.42233037072213, 0.956339100654794, 
    5.68982662883706, 2.8189887994052, 5.28333523725378, -2.15455097416025,
  -9.11738292082699, -7.65290582112484, -0.271904391569432, 11.2325459788246, 
    1.51637228367027, -1.32881403833835, 2.22954506335454, -8.46592050769422, 
    0.400129652303432, 4.49353871319253, -4.28290490508767, 
    -2.55692344457882, 2.84501739136846, 8.89256569445797, 5.64104336225571, 
    -11.8954098259313, 1.06374037794511, 7.98911186743826, 8.03469018056542, 
    5.82355103744084, -5.17114284457893, -10.7355828528363, 
    -5.72534094057754, -2.33292670670801, 5.81058656303432, 11.8129856383325, 
    4.24883441201218, -6.82372992657744, -7.55277515986734, 
    -6.37596958769715, 1.12391460041977, 12.2776681256866, 7.54737772655331, 
    -6.00587063510384, -3.58411629177168, -3.10256302403837, 
    -7.53267058732873, -3.99540411170554, 3.76074484956272, 7.38250135993267, 
    3.47114877746848, -3.12275338709991, -5.71842534290698, 
    -0.166564014173535, 7.76735404703243, 8.42861720475397, 
    -5.31910957727861, -3.90264208673532, -2.79921564854511, 
    -7.78344519525623, -1.40425024956342, 7.31917626172761, 10.3863768398576, 
    -1.1004095363927, -12.0658143210842, -9.29349746999864, 3.58410175174658, 
    8.43128545219046, 7.20018407749626, -1.77413855018538,
  -7.70416460690991, -12.216433436989, 2.80985212971745, 15.0399649808913, 
    -0.693130246992926, -3.11590526763342, -2.15297587392617, 
    -2.80923242442632, -1.02430864428147, 1.27277513107891, 
    -1.16043479024954, -1.73626993656586, 5.91384615137578, 4.14119617374593, 
    1.70337514323, -1.77338693533411, -4.74219830773553, 6.07256143190931, 
    7.70424098064429, 2.28686687381677, -6.16949888848091, -9.54856855594024, 
    0.647220836018436, -0.3652975069709, 7.86840515407462, 15.4336231772184, 
    0.00504005082462495, -16.2085145987437, -12.5298862323092, 
    -4.31307819225679, 2.10418194535244, 12.8281794942926, 7.03065788476951, 
    -2.55875093494489, -4.00155372865643, -2.83163141778234, 
    -5.49334771973057, -2.3995118722459, 8.08552923368994, 6.70528127801436, 
    0.200022175070057, -5.32196876478505, -8.94512247381647, 
    -2.01901287533932, 11.1421509608511, 7.63552222744724, -8.30296588419151, 
    -2.01869244495045, 2.09898243251367, -4.39350176247703, 
    -1.71219506167834, 10.8257239766189, 8.29217066147006, -9.01545851592804, 
    -11.9245680685904, -8.73975753479964, 1.70362637515442, 14.1445093309466, 
    5.9889774675621, -3.99189959993752,
  -8.57276356097765, -9.45736736210293, 7.81302522282355, 9.56181363103288, 
    -0.392743694700267, -1.02750403219893, -10.0247024373203, 
    2.24207608795533, 4.4678117015484, 4.81110750983455, 0.814352903516753, 
    -2.40913927550166, 0.485295332576845, -2.57392958208255, 
    2.93144625024061, 0.977069526106712, -0.931558803196134, 
    11.9948731821387, 1.24154119309962, -3.79176589000464, -5.40635397687231, 
    -10.075098014333, 4.34375912990917, 4.90119474665649, 17.2024203700402, 
    7.71782443793819, -6.99041194782664, -17.8657348218111, 
    -13.6684068426598, -6.54413347274936, 7.14594081344092, 12.170643725549, 
    11.1716587081072, 0.0703788641509251, -4.31911752753835, 
    -3.79101884644302, -8.58718762181683, 3.25636280633082, 11.4761177881707, 
    4.65737143784135, -4.99287077471133, -8.58750654903026, 
    -9.47088533346861, 2.69740577854979, 12.4191602921321, 5.09374133469082, 
    -5.15342686762559, 0.578648614061451, -1.51640246511003, 
    -8.65149339967534, 7.9505123068055, 13.0415908699037, -0.328042344621423, 
    -7.9045127712093, -14.7128515314235, -6.09133749679383, 6.73069521379461, 
    15.9820350295544, 2.54933213872497, -9.11684698744472,
  -6.557674857471, -4.99777613286406, 7.86110457869674, 4.27444757316523, 
    -1.54858514928076, 3.56087783693785, -3.53581386134635, 
    0.883854914276704, 11.9604898300001, 4.15282210998835, -9.94051511955535, 
    -3.70894480407894, -2.07155874829024, -4.24541304851069, 
    3.62404932432297, 5.34266221715543, 9.12572106693373, 9.71122676204647, 
    -19.8718866569807, -10.9136216573752, 1.05211929045366, 
    -8.23245876923841, 4.89570610928825, 17.0638872756732, 13.6871240455805, 
    -4.69531620298609, -8.86898432924165, -12.60602749412, -1.92372172769228, 
    -2.32280313663725, 7.78887635432807, 12.8623471123924, 4.27227173645771, 
    -7.94612885366732, -3.03462737688061, 1.16490822614018, 
    -6.07720302392871, 4.53657085647931, 10.3866137731415, 4.13549402442951, 
    -6.63132094443005, -7.97843814906736, -3.97402866336306, 
    5.53905396783705, 7.81420976491656, -0.334615439704745, 
    -3.87251082066366, 3.43435367009047, -1.75734999893511, 
    -6.75180031155541, 13.5776939972718, 9.07795621887, -6.78760908705956, 
    -8.57340534464279, -9.18245179653448, -2.45287909906774, 
    12.4877008976149, 8.6780841596874, -0.545130030600607, -9.67605691878583,
  0.428697019283364, 0.162110449312061, 4.61367187492671, 4.65290581062502, 
    -2.13734969521743, 1.78815480694515, -0.952407749484849, 
    2.02920032229513, -0.130442909990905, -2.57492051424268, 
    -5.0338045968391, -1.63172707803215, 1.86280708596898, 1.75665306519085, 
    -1.21384994347769, 6.27353333679747, 5.60763463262769, -1.86737242990829, 
    -14.3842788470861, -12.0725526190426, 4.20156508083256, 3.70539303012091, 
    -4.08950542630175, 11.5022396985326, -0.382844736294405, 
    -14.8970610515027, -4.54725888496107, -5.73481909301279, 
    3.23145502829483, 2.81084419254771, 2.76250297765794, 1.073477571659, 
    -4.19668030735262, -7.23290605314147, -0.255656295251244, 
    2.47474026708781, 0.150961059927619, 2.15303205377035, 6.74568287881894, 
    -2.37412368112439, -4.22791296698959, -4.85857272957967, 
    2.91541873693149, 4.71550447731361, 0.199424676697876, 
    -0.155019389537246, 0.661985572396976, 2.60882198543133, 
    -2.99901508695837, -1.37023596581355, 8.76125462668412, 0.28370099289433, 
    -4.40415685984948, -3.35616007958792, 0.0465664493073245, 
    0.602141423769629, 9.00509444132056, 1.82053765115031, 3.14232843928484, 
    -13.4590504693013,
  3.16721438257025, 2.45914000268421, 3.07127535460042, 4.28694331364815, 
    -3.73077166111769, -9.12300823438069, 3.80077319863674, 
    -6.22675424152113, -15.8919420199547, -7.15219614167868, 
    -1.45460375511084, -0.966115634597579, -1.38225862132511, 
    3.48968532011291, -0.0180975338676081, -2.84414129372328, 
    -8.38434119763106, -9.30816857023779, 4.37393383438865, 
    -5.87103222822478, -2.40481253923378, 1.98621741874079, 
    -2.30141391578128, -1.25256666580151, -10.9224153589402, 
    -8.19247810820583, 0.367454861549341, -3.17499905517713, 
    6.92705242796771, 3.29892430981193, -1.57941020921092, -5.37094256035131, 
    -2.37826806679104, 0.0203527431780853, -1.14720896932384, 
    0.613771647123486, -1.20215598016478, -3.58903927345103, 
    0.918814871690043, -5.52949387914319, -0.00157872760581736, 
    -2.13424800539391, -0.5771236037236, 0.939921747606176, 
    -1.58570527827339, 1.14051372248666, 2.48873825448525, -1.01779376981973, 
    -0.602280347879546, 2.44112446972738, -0.623062963716743, 
    -3.60891829630381, -2.87050522953171, 0.291966111727008, 
    -1.50363316965022, -1.94351541901623, 1.66457596077608, 1.58467589360063, 
    6.87325106786729, -13.0403732283104,
  -4.48746964813653, 0.673810952931338, 0.560036240705279, -6.27679756224961, 
    -7.6147574156456, -3.53029491806976, 9.49682404216376, 13.9744550067244, 
    6.85880056328818, -6.83143920901088, -3.58934756994436, 
    -4.46656909946334, -5.20379726811559, -2.56093955624769, 
    -4.49483767095667, -7.29827277492954, -1.80697580757135, 
    -6.91737119221027, -0.081825627555727, -0.413419981335449, 
    -3.83813693621137, -4.02089697131101, -4.50148882271511, 
    -5.25199573930569, -2.89603220656091, -2.81970898374285, 
    1.99623147554448, 5.25198321424315, 7.21228029451517, 0.487476956130244, 
    0.130675839027179, 1.18697702967725, 1.85862872100053, 2.45088816351001, 
    0.04436246401838, -1.47838063677074, -7.06772580815099, -3.1008607209102, 
    -0.528440142049448, -0.117442805727322, 4.95107009017869, 
    4.67717449433991, -2.27171680077119, -5.28565277827859, 
    -2.49837560618229, -1.57139159462231, -2.38955328421359, 
    -7.06812952042235, -3.70276953445095, -0.642285164498669, 
    -2.50257548784796, -2.6949268166284, -0.683913981888391, 
    1.07435627008605, -0.185776585190833, -2.13061481533958, 
    0.63082750414041, 5.09518805189368, 10.2416853782214, -11.2588164439931,
  -7.81296561020791, 2.90247120212154, -0.882677276529885, -5.81115205626069, 
    2.1279787848951, 8.48632733878698, 2.42029523358788, -0.678148767763235, 
    1.45869633299285, 2.23883449069046, 5.34651506610868, -0.689495343895975, 
    -4.73164021697232, -1.18294962933503, -1.2133098733724, 
    -0.946392108827449, -0.881956497990181, 1.78799770710359, 
    -3.34130995685342, 4.42286220625986, -1.82861189674206, 
    -4.59876066510919, 4.94456095417844, -1.6220095805761, 0.659343835937158, 
    -4.01265505285943, 0.225727475996733, 7.31008435046266, 3.16125556221843, 
    -4.66591038067894, -4.68431579863835, 1.72283669820172, 
    0.330801631137667, 0.887452348740709, -0.272517230679344, 
    2.89623320541271, -1.93942943948545, 0.339422544073163, 
    0.206213005948806, -1.88814743943639, 3.83005851508609, 6.70679003099354, 
    2.75467069592633, -3.33187771617634, -4.50048016783656, 
    -2.14863506405526, -0.249179093585259, -1.72021361750598, 
    -0.965431790961505, 0.800325764920091, -0.470131505895786, 
    0.293653142375204, 3.11030258541391, 0.737103346136859, 1.51268627004726, 
    2.16022126987998, 0.759347311283642, -5.22006332523044, 2.127391678384, 
    -6.51623464922527,
  -7.98249711323363, 5.6855577182097, 6.17446927482839, -3.2867126526418, 
    -0.773085269514311, 4.48600938572832, 4.63123583382354, 
    -4.77481437136627, -5.9614801008594, -3.28589704454332, 4.31172860598682, 
    2.88548995178314, -6.43692772637318, -0.117075271874229, 
    2.94155676555515, 3.59599231864736, 1.25353775077772, 0.631810185073815, 
    -2.97720338739031, 2.93324644410624, 0.110535721003994, 
    -4.59703825182763, -0.578434048032815, 2.74029608141969, 
    1.78394758827251, -2.44457525896306, -0.804625357082149, 
    1.60528730569908, 2.60035916177475, 0.777046144155799, -5.48592940700772, 
    0.820251113819819, 9.20277287668588, -0.516806474493745, 
    -1.62937651024268, 1.88364688166193, -1.36466598276271, 
    -1.80642044242685, -1.21651135893278, -3.37946679878865, 
    -0.209683425629947, 3.75465679087016, 0.26315240125893, 1.70389615927253, 
    0.448063191834391, -4.1260136750619, -2.23970382073509, 
    0.900502689631275, 2.31560205491886, 2.27234689955942, 0.157383867535861, 
    -1.31585924743101, 0.388825794754611, 0.835815166387059, 
    0.849015596602855, 2.10551094130876, 1.60281892360263, -5.00100501094072, 
    4.51708311314784, 6.65210847872975,
  -5.60636566097145, -1.95290673210387, -0.41431840530862, 1.17471721775312, 
    0.997535856870666, 1.72035913649439, 3.36264551048685, -5.52850319372668, 
    -9.51165302992513, -5.87707525741903, 7.42926725597569, 10.3907189040548, 
    -4.99528982817424, -4.17724452521918, 1.4917585922236, 3.28848721051765, 
    3.25929294856843, 0.422065220611914, -7.29486256958049, 
    -0.271083293685491, 5.8925565578496, -1.18888253145977, 
    -5.10116361707786, 2.09195010552949, 2.36078668093227, 1.10585339533913, 
    1.15492619288787, -3.62022203350447, -2.42357883319197, -2.0676795067951, 
    -4.26927434464135, -5.20395318304537, 12.667791991635, 5.43162017624997, 
    2.04583122761712, 5.9084918560911, -1.92006800402141, -8.34829888593225, 
    -9.67512724503818, -5.1518227096589, 2.34939414756906, 5.17579277991345, 
    3.42869147041571, 1.35857935243278, -1.54939433402842, -4.14289918758051, 
    -5.78798997375078, -0.468314491320714, 6.27281691111773, 
    1.06775766910397, 0.751080654796705, 3.91101821367606, 1.00791285818567, 
    0.718457962085513, 0.944138548065155, -3.92002531122885, 
    -5.63282013370214, -7.2387604203051, 7.47227189433626, 9.55737378313397,
  6.37340482296209, -4.25437292150951, -11.4405019597905, 1.91290699140817, 
    6.46244488447909, 6.67321064427775, 5.70395687103351, -3.98014081014702, 
    -15.5505757521099, -13.5628009064885, 5.31695312730169, 14.913739061642, 
    3.299282178495, 1.18398543226152, -2.53805467350378, -4.21767588232427, 
    -0.594727071187891, 3.46337668820907, -4.21070648203329, 
    2.22295681601602, 6.02662231459245, -1.24362779336336, -7.21668056904831, 
    0.509176112529549, 6.179920580652, -3.24986325399369, 0.214991566561585, 
    -2.6568638926246, -0.335243603335823, -1.82392351182923, 
    -1.14402029207656, -9.57603892486308, 0.35660590711107, 10.9359655362566, 
    10.346525532331, 7.25412265340011, -1.62710484455223, -6.80171892668581, 
    -10.2877673959668, -9.21935322533397, 1.93272491497735, 6.86731676891298, 
    7.48693893613538, 2.98826780444151, -3.51583127588498, 0.340048437474744, 
    -6.00987717509882, -7.37383478620988, 4.85124520867778, 4.06743568127434, 
    -2.4150500527006, 5.39272190833589, 5.52442734021237, 0.811905708841746, 
    1.12612617965964, -4.32298217216285, -10.5764954347869, 
    -13.5496834867988, 8.27589185533922, 8.45676441916919,
  7.32388536238287, 1.20678134617161, -7.04173318776476, -3.2244802233787, 
    7.17801463964314, 13.4237001956207, 4.52354102397763, -5.2418657917278, 
    -12.9853082093442, -17.8416454880167, -2.43394074185926, 
    13.0175129229154, 14.3986987959845, 10.3454885673128, -0.81083837412439, 
    -12.1270462720697, -9.5752281566372, 4.36929167057286, 5.23049564717336, 
    4.27097999637204, 6.13127721420188, -2.80247875027841, -12.4767824311713, 
    -3.31383460547431, 10.0847568798753, -2.71557585516343, 
    -3.40727776210097, -4.10076310267965, 1.48688460874202, 2.59972033519363, 
    1.15845782190641, -5.78491912159032, -8.14929468092898, 6.58502933430297, 
    11.7444584643421, 3.94967393974917, 2.02088166432375, -3.2752390809731, 
    -8.52051082430924, -7.31290188088548, -0.250384932649747, 
    4.46579077220162, 7.29597572601136, 6.43928458956351, 0.250385950724468, 
    -0.884219204912045, -1.87734850656334, -6.6126786522906, 
    0.340386427471978, 5.99883040042845, -4.51957957670316, 
    -1.78854863051666, 4.03330628456276, 1.35421711645162, 
    -0.691987580118169, -3.2148485493648, -9.90661721965211, 
    -15.5233936687351, 3.50748062097176, 14.9139853384621,
  3.35370772379923, -0.436007315227718, -4.31295624707837, -3.25487267770222, 
    7.22578055429955, 9.45983442616566, 4.65446493572715, -2.48451176876316, 
    -7.55481380010744, -14.6440152801561, -5.56219535100459, 
    12.6316656444003, 14.9949989522221, 11.4145671851398, 1.03036912969764, 
    -13.7070581473627, -13.6482545480465, 1.17100164282358, 11.2156999039945, 
    5.48240270139792, 7.62554119541962, -2.57446120698904, -15.7838806886711, 
    -7.76967235441979, 4.29719905926223, 7.22287099433177, 
    -0.680709431028884, -4.64670356823663, 1.91967909722877, 
    0.956712502462265, -1.99500447865809, -4.23913142327165, 
    -7.17765129088907, 1.1835380749374, 9.12098788595133, 7.45630001821964, 
    9.23544724545786, -2.07535822517175, -11.3111108839787, 
    -5.70501210113238, -0.85822057711862, 1.45616606582751, 6.26099705594497, 
    7.36204182833016, 5.19137325602418, -4.00690430093368, -2.05718538675949, 
    -1.73690476083204, -3.33728703430475, 0.243636713230154, 
    -1.05427438398847, -6.78083952268735, 4.4193175104219, 5.03612698529691, 
    -5.32457285844964, 2.35663401323983, -3.97643051723961, 
    -9.13563271326892, -3.13106838064091, 8.19074080496643,
  -3.52618504934905, -2.16902833081459, -4.01929390430989, -1.82784490151113, 
    6.29683759553826, 8.42902260448237, 9.71861367568625, -0.836018577839125, 
    -8.46310563140223, -7.80911312685515, -2.95910686127231, 
    10.9174044372576, 9.13964460581758, 7.38184591714888, 2.18489006732281, 
    -6.14787994936725, -11.3188551728392, -4.76940320376242, 
    4.94985687652383, 7.23734919811433, 7.4143707502386, -5.26993118117348, 
    -13.7660232636594, -8.41091109973081, 5.14028614321777, 11.3354711734631, 
    2.28951158218355, 2.41104017599606, 0.937510491623179, -3.73444903673135, 
    -6.06045649855985, -5.24412020732991, -4.81828907419228, 
    0.136044299144582, 8.15003227085215, 10.4626841143822, 5.9090739922667, 
    -3.60480292296233, -6.63882282893256, -3.45957306711093, 
    -1.58504072616416, -4.06141121565319, 4.14982206839215, 10.6328988750231, 
    7.32552699322925, -1.52540701363035, -4.80679595158863, 
    -6.10527314616335, -9.0029982797637, -4.4079895203098, 
    0.0267430085920801, -5.20659022614418, 5.02370087730969, 
    8.24712582896884, 4.16825245244976, 10.0335555545801, 2.68923064282929, 
    -5.33837324553299, -8.06120383759247, -6.64705950759267,
  -3.76033999440072, -1.5061053871331, -0.875008415912433, 
    -0.273886985777993, 5.64026883575697, 8.21021812951534, 3.03658534827731, 
    -4.67219352500983, -4.73223743557964, -0.319753216033639, 
    2.41866047527421, 6.67324802995061, 5.09814448483826, 2.77121921027374, 
    1.40849004271497, -3.45163621144802, -6.73716442532236, 
    -4.23285067370113, -1.18004439744283, 1.11467443592794, 
    -2.06595995421168, -2.70012063616527, -4.4312448636504, 
    -2.27149563885366, 8.68037671634194, 7.28395428565866, 5.39236912526916, 
    5.04036826419809, -1.94410880129204, -1.34919888827541, 
    -4.36918117257066, -3.63088131563066, -1.65108194884095, 
    1.82500384196941, 5.12058718571017, 3.70937005678087, -2.47494793683767, 
    -5.80768180193559, -2.83912915511497, -2.87841488634851, 
    -2.63412561358378, -0.728677072132407, 6.2501447939749, 11.9098341313161, 
    3.74613395292811, -2.10824769482544, -10.5899880837548, 
    -11.0228970406589, -5.23986812734299, -0.668985577540584, 
    -2.36060887275901, -2.80723162908683, 2.9358295258343, 10.2072254743599, 
    12.4094655675659, 8.81649625635197, 3.98679178756905, -4.81735923489115, 
    -8.50642377543741, -8.33552469573159,
  3.46010576933196, 1.98472716300119, 0.144126911805685, 0.413717507057144, 
    2.28187487118654, -1.08687189287792, -5.53417010282207, 
    -2.18692418895672, 1.29320414429253, 3.31116421820248, 3.82282504890427, 
    4.19239403263981, 1.79950239673395, -0.738366857409461, 
    -3.47382503542859, -8.63582988475897, -6.12196045522602, 
    -1.25582120024605, -0.147566932465088, -2.03970415024765, 
    -3.17751939973333, 3.36955137686633, 6.25455057444732, 3.03600539289544, 
    3.67194072254901, 3.38087592943919, 4.36038785461945, 0.653125200771063, 
    -0.866193738772242, 1.10567941011363, 0.493633992601276, 
    1.91669681106975, 2.26036215248054, -0.195218415230241, 
    -0.694930706203083, -3.6200746144705, -9.77642980769207, 
    -10.3745014377871, -0.431334776844398, 1.44190364875491, 
    0.742881891509471, 9.85748059261272, 9.91364870743818, 4.66392208707668, 
    -1.59778224342172, -3.77209017871256, -9.62068383401656, 
    -3.23266532181666, 2.66993333387324, -3.54829222806448, -5.590816277327, 
    0.557841954434223, 2.36227029513758, 4.75707257670343, 4.28119994078308, 
    5.17227616787274, 5.88430036431191, -2.15930007889133, -8.2616189734424, 
    -4.81795799972345,
  5.69487156514583, 4.83509871013264, 2.67676001569675, 2.6604686371936, 
    0.0376769984782261, -5.30398404396381, -7.30084566482412, 
    -3.5524713339892, 2.60756871045991, 5.08396607455996, 3.65431450005428, 
    2.93341762368375, 1.01040635841921, -2.82530184073546, -6.62804060467268, 
    -9.62683807826158, -6.80782806364621, -0.499699321509275, 
    1.92548783445213, 3.34298929443557, 5.06706327625183, 5.55145573569282, 
    4.85189488996548, 3.29737515246165, 2.46324141028511, 1.38941919506838, 
    -1.32959201822592, -3.38202043687892, -2.28086674074798, 
    0.184882954421022, 1.87519450011689, 2.81193738803843, 1.64560528961166, 
    -1.1752545686528, -1.08000975638359, -2.1793896402226, -11.6249399076043, 
    -13.8100473657133, 1.61399395709329, 10.1564205691644, 10.3416731498948, 
    13.4237495277559, 8.14505240914536, -0.380399023309346, 
    -3.66708144585177, -6.62962556999055, -5.17630359922469, 
    2.79849932398424, 3.82143507182741, -3.59287566026057, -4.91233682785022, 
    -2.65144297558006, -2.65935221353691, -0.436504960318242, 
    1.39283225833009, 1.61166923731424, 2.14001829155946, -0.999680426956709, 
    -5.28489644265707, -0.485822982075761,
  4.1222047231172, 5.28477047774026, 5.66142644061536, 5.04840984397373, 
    1.60816643529478, -4.0435216541702, -7.55040173636002, -5.85189221127621, 
    -1.31727199173488, 2.16398765406736, 3.53566127512366, 3.84116187921061, 
    2.99189433546016, -0.427226993056498, -5.85715190955919, 
    -9.13575188074674, -6.61450621362611, -0.232516861574285, 
    4.74549341438235, 6.34105635588872, 6.03377152276128, 5.49045293173418, 
    5.21082516642324, 5.02038975314702, 3.93990640349525, 0.698913975670693, 
    -4.09354859466521, -7.54363218414868, -7.357600074085, -4.2505176950516, 
    -1.40057636783171, -1.26218270635256, -2.18082869332949, 
    -0.347421989066947, 3.3171076071027, 2.50249813722399, -4.06236052701384, 
    -7.53831895506225, -1.52411661843688, 8.44611820701893, 13.6485134813143, 
    12.9904703781517, 8.07088730728908, 1.07702769852791, -4.55053085818726, 
    -6.79615692997472, -5.78767254848474, -2.12916702815351, 
    2.00942765032373, 2.35507961207257, -2.19999849196691, -5.76988221500578, 
    -3.7958217090907, 0.08022398994094, 0.812814808855009, -1.30010190097818, 
    -3.31584683357646, -3.60297380506087, -1.87976900553147, 1.29498726598671,
  1.56652666246808, 3.72883778803596, 4.64368983475958, 4.59171069087624, 
    3.39133574713565, 0.832900819363069, -2.51031533300633, 
    -5.08903355915924, -5.42968093485231, -3.3955799233104, 
    -0.209615104834303, 2.30591864475835, 2.71932800156717, 0.84350037912604, 
    -1.84746962933263, -3.09074111084377, -1.58765185880977, 
    1.88132315642246, 5.00224516970883, 6.13692871178138, 5.73624676849814, 
    5.28973361503501, 5.47442501032747, 5.41080864617312, 3.55367952287765, 
    -0.595227853332462, -5.62947143364704, -9.06493989032436, 
    -9.34231287105115, -7.17476220902215, -4.61489610882768, 
    -2.84552667211528, -1.22888933800425, 1.20239214695046, 3.80061787183364, 
    4.65335966895642, 2.83195528040741, -0.10822015822434, -1.44789742561664, 
    0.414546499232002, 3.98574357971959, 5.98987779690308, 4.71177475163461, 
    1.20652730165961, -2.04144686126129, -3.25975898371934, 
    -2.47001285560908, -0.953221281263259, 0.133003458813475, 
    0.492314245869405, 0.363418522621442, 0.283710801036074, 
    0.824866890849863, 1.49012579101554, 0.833507179564416, 
    -1.73683494827992, -4.90402457171277, -6.4129811570098, -5.0988074157481, 
    -1.80257396564648,
  -1.19164938724995, 0.721901672744847, 2.40453729838361, 3.32701220679117, 
    3.19064814851777, 1.99521294173428, 0.0925185670140736, 
    -1.93971831517063, -3.47028120232455, -3.98395717746849, 
    -3.39170104627575, -2.07632031241056, -0.621314704905249, 
    0.529664800153096, 1.21004502674941, 1.55406037802456, 1.82114226983609, 
    2.20298383105618, 2.74247603767845, 3.2985959085139, 3.5888741357536, 
    3.37881466311094, 2.56708673370967, 1.2379620329563, -0.355532876586324, 
    -1.8934682648665, -3.11595461547876, -3.87887229826166, 
    -4.08364423064782, -3.67152682856935, -2.665202113826, -1.22470632622171, 
    0.340322726433255, 1.66323958384965, 2.43925490088416, 2.47888712633158, 
    1.81348024602221, 0.743163031477657, -0.37974143945842, 
    -1.23630620879771, -1.55892791238778, -1.34558291340485, 
    -0.865372320565576, -0.428937563336063, -0.210032990304099, 
    -0.20049494221209, -0.281685728260665, -0.30710073441302, 
    -0.109646064996155, 0.385167754874833, 1.12871893353323, 
    1.96330201146126, 2.50317184033622, 2.38121981776311, 1.48555889468464, 
    -0.00422016803691948, -1.64583230961146, -2.8976722736013, 
    -3.32014162439873, -2.70553047097173,
  1.04669758997801, 0.794160123683808, 0.505645187985983, 0.201406169379881, 
    -0.10388113124984, -0.383996836746396, -0.619710341591498, 
    -0.79682682632713, -0.906184389043195, -0.956346601329453, 
    -0.943441193333188, -0.856601081677478, -0.697335449760635, 
    -0.490503970713728, -0.271822209081792, -0.0759991798386218, 
    0.0700038561385714, 0.159369170870569, 0.199655177487297, 
    0.204221764832765, 0.197030356571436, 0.199004399573465, 
    0.229343447238863, 0.301901863595431, 0.412859657845558, 
    0.546228888668376, 0.677155126369616, 0.769857396408008, 
    0.782456109821789, 0.686993196104942, 0.478458101319248, 
    0.184362918159544, -0.142685173207811, -0.444055787488956, 
    -0.67141653562549, -0.788386135011583, -0.785611720840356, 
    -0.678736792167859, -0.496670144257595, -0.286980290641832, 
    -0.110313650256435, -0.00350355559808129, 0.0291051444074427, 
    -0.00530076349847017, -0.104274725914863, -0.255847651735748, 
    -0.426391756396998, -0.568597559266403, -0.645768083104534, 
    -0.623392050305921, -0.48845724456051, -0.273793219237222, 
    0.00590522877255062, 0.328068443958522, 0.644343394194879, 
    0.914563213607585, 1.12482866220698, 1.26373412844523, 1.3049608236185, 
    1.22923951093239,
  -1.51849676165507, -3.11547150905098, -4.65619291948144, -6.03221882994714, 
    -7.12237340362014, -7.80705888961559, -8.04030204702497, 
    -7.85142694980618, -7.27440802600898, -6.35625163948213, 
    -5.17054418951559, -3.82465734574347, -2.44374691850556, 
    -1.16219532480197, -0.0956793493634283, 0.681793093892173, 
    1.14254311353711, 1.27694787859117, 1.14030660374694, 0.850331895497799, 
    0.531359225008883, 0.27900301589152, 0.143269009876858, 
    0.154072564554462, 0.323899508293048, 0.666087581157377, 
    1.18078795625686, 1.82140267350768, 2.47951738941899, 3.08536462461099, 
    3.58354700281421, 3.86730004765823, 3.87879832076927, 3.63448240585174, 
    3.16570898243641, 2.51394591747897, 1.73459965240189, 0.895818549712964, 
    0.0616652942030312, -0.702929165471488, -1.31028383835471, 
    -1.69089516424808, -1.81370591677008, -1.67196041116612, 
    -1.2765623164168, -0.645734760826277, 0.196246308552834, 
    1.19287697393656, 2.25461969658595, 3.27571571409681, 4.16687057301039, 
    4.85179410297368, 5.27128614101851, 5.39122351574581, 5.18931818815115, 
    4.6757755966203, 3.87525659599247, 2.81539475417909, 1.52662445312183, 
    0.0549750544994309,
  -3.78422067140422, -4.74453675483518, -5.01509065478164, -4.72793568105526, 
    -4.24040267119676, -3.96799032804496, -3.96795323424093, 
    -3.8813298140544, -3.37228976702846, -2.46736988729493, 
    -1.58289034820019, -1.1388254021857, -1.23694896674887, 
    -1.63345486374996, -1.9852511915721, -2.02850417022136, 
    -1.64680522243924, -0.777912067148072, 0.524898623703138, 
    1.65679045016579, 1.88600808203864, 1.28030091699281, 0.529527625676043, 
    0.25752385717849, 0.737595277197873, 1.78124518527235, 2.89180575873725, 
    3.58496755801325, 3.72273121241825, 3.38399116119288, 2.85567764558518, 
    2.650947870314, 3.00585805797317, 3.68162402519205, 4.19917851265254, 
    4.06353009757623, 2.98163171175483, 1.00745735666757, -1.45290075681696, 
    -3.83947744081704, -5.66339238752366, -6.49088312205427, 
    -6.00825092614575, -4.244640378721, -1.67330865313973, 0.978103855172097, 
    3.05051188989525, 4.16786725517313, 4.28658597584517, 3.69851423352585, 
    2.86791074044746, 2.24344237793507, 2.07343108319904, 2.31116800246955, 
    2.71040384299842, 2.88630347088631, 2.46435736805335, 1.28024584232545, 
    -0.446479997403882, -2.26138665071869,
  -3.49067246720699, -1.72353001032833, -0.25544886354391, 
    -0.731433540708513, -2.18790812729448, -1.69485095110461, 
    1.7802405585819, 5.46577733625741, 5.70620958613267, 1.85586865356734, 
    -3.09529164445295, -5.6874211002656, -5.54825448933785, -4.6326895312981, 
    -3.76633433876462, -1.58117561763939, 2.72233285677061, 6.75199998759674, 
    7.17248808900553, 3.96302436798873, 0.449228220077085, -1.0793876714026, 
    -1.35175391135915, -1.3731748026473, -0.785121284086486, 
    1.03743321218978, 3.33751419665066, 3.95491711641635, 1.47959903907202, 
    -2.23852100475069, -3.6491964217064, -1.28375643396411, 2.73764212297939, 
    5.1055100101957, 4.48912653076513, 2.22429704724748, 0.537433973191825, 
    0.232194306066206, -0.335787624992167, -3.04560310363827, 
    -6.9286277714924, -9.18289751600657, -8.08206828655629, 
    -4.07112768352587, 0.745184520946308, 4.03741174764679, 4.73187817201123, 
    3.55675601809508, 2.33739352232661, 2.17750726473444, 2.48650128601391, 
    2.16448643067205, 1.19149948150773, 0.352516175746372, 0.112693163662408, 
    0.246718286041109, -0.0140319100509878, -1.0010174077069, 
    -2.49604192176264, -3.73971087236192,
  -0.51609209267463, 5.0188456977561, 3.11921853288323, -1.9269653841799, 
    -1.92760551151299, 2.95676053683417, 7.99580638980341, 10.4967767503193, 
    7.85093344623615, -1.06716930681077, -10.6400900749973, 
    -14.3166201865901, -12.0031285764181, -7.23787619678641, 
    -1.2197492352209, 6.85935925193618, 12.616001117864, 10.5314293980157, 
    2.98152562550675, -2.89991432016583, -4.29595723828742, 
    -2.50122906374567, -1.44191223031762, -2.65394367311781, 
    -1.29647749276374, 4.06177861773806, 4.63941864868982, -3.50747844829411, 
    -8.24240269195479, -2.82006514062566, 2.15294002764446, 
    0.718299705181413, 0.168506629796196, 2.68649764817441, 2.23191144978471, 
    -0.134413634174865, 1.85847149455194, 4.6619126540618, 1.10558658700484, 
    -5.15444572776844, -7.45600922503071, -6.6967203526606, 
    -5.11099976272911, -0.855366936131699, 4.77758367016403, 
    6.19579691763407, 3.47447926616941, 3.09948295734009, 6.14056369032152, 
    5.77358346676076, -0.715453773662691, -5.68381648516631, 
    -3.45707140594409, 0.0317408438029192, -0.389691125549341, 
    -0.406405937464866, 2.3702559117397, 1.69062377969896, -4.06748074747219, 
    -6.20048515777767,
  -0.727198922140049, 4.58951318846778, 1.2579031903161, -1.68265271297541, 
    3.04339125404088, 6.52371768410791, 10.4375661444122, 14.7379260153853, 
    8.52841942950895, -2.87093525514555, -9.91287192312964, 
    -17.6817930346809, -17.6112180600384, -6.46698492896704, 
    4.52783525118004, 12.6325088184037, 12.1254785752016, 0.336286246325499, 
    -5.0981939398642, -5.2501949547899, -10.290189224171, -9.8722087160169, 
    -0.161615154180316, 1.62136953556754, 2.24594267001806, 7.85269537607853, 
    0.972067488421716, -7.96648529294019, -1.89787323324448, 
    4.05175995531969, 2.17682207829325, -0.214316829892458, 
    -1.22167147052339, -1.8885881290963, -1.56879110344558, 3.19484619215416, 
    7.28138397791891, 2.41625789586172, -3.27186730542706, -5.50091481496032, 
    -6.46790440176736, -3.59176883471494, 0.428672048927343, 
    3.75899193510771, 6.35875844916063, 4.41714338912989, 1.4241418900752, 
    4.02298289624396, 8.97265099103509, 5.21150607979045, -7.60546789697432, 
    -13.1091729529816, -6.53097906052832, 0.118876259110078, 
    2.18759211138216, 5.17157165609092, 4.38048175617081, -2.4589508885907, 
    -5.44775534574643, -4.47806142807403,
  -4.00169175737498, 1.65330935520367, 1.87644196719388, 2.90939688765283, 
    4.64727486698554, 3.98944239417128, 4.81343237809645, 13.9307716168788, 
    12.7284751585637, 2.30332306066965, -4.98146321887423, -14.2657634416532, 
    -15.7026725570424, -13.8306540687242, 9.87478042751978, 8.99381681731165, 
    7.32314244370054, -2.35327784581991, 1.70793648144674, -5.11287430036598, 
    -12.42490119655, -16.7763038846902, -2.70848621999055, 
    -0.470005792502501, 3.14420050946554, 5.58124594940193, 
    -0.79330964325534, 2.32154893826561, 11.5456430386462, 3.40717790352556, 
    -6.97839193537174, -8.10996484531872, -1.555227246292, 
    -0.594332171672018, 1.62536678197759, 8.34097066099706, 6.96138695261571, 
    -1.01446723056499, -5.54973937178085, -5.57172849881761, 
    -3.56306768008374, -0.778184104359317, 3.69674139009717, 
    5.02349066976972, 5.25596237384165, 2.92353766188484, 0.671192997992288, 
    0.796939883494499, 3.62791895767324, 3.89884610901139, -2.29324952182627, 
    -9.62701836056679, -11.1988132198215, 2.49934364604246, 8.12790350114146, 
    10.7194044528453, 3.73381482612478, -4.05172130523607, -8.18552789919338, 
    -2.64215721502314,
  -3.43890528375752, -5.55980791308479, 0.18854311055082, 1.14423830598707, 
    3.10714968447477, 1.60333444665101, 0.87114650367056, 6.4630219409273, 
    9.57991923760688, 5.64113533846377, 1.30174650723193, -13.9391545463248, 
    -1.60990973127999, -12.628632509261, -1.02742399893058, 6.81477508419756, 
    6.35583599610565, 5.97128373588611, 10.2872564380357, -4.79314678622225, 
    -9.85277816982963, -18.2929586522769, -9.91859616975855, 
    -5.23055402994721, 0.184241408554302, 3.20029149622043, 5.42180866178466, 
    11.4191600396686, 10.383314941392, 1.52402062614901, -6.68814777962105, 
    -9.48179780947438, -3.33437616492601, 2.17469914067477, 3.85297534200923, 
    5.4207939998321, 3.90390532899506, 0.420687107890335, 0.256287233117797, 
    -1.38961546378411, -3.59354705454108, -2.44592608622463, 
    2.35290854591532, 4.95624066645827, 6.16212099924883, 4.09276323935669, 
    0.611778475229818, -3.49353608523963, -5.48361502837325, 
    1.98065698925148, 3.6616208164058, 1.34250606617808, -9.51081388028843, 
    -6.17855394183682, 8.61410941905768, 8.55101908702007, 4.76162383235393, 
    -1.29752089941678, -2.0041499995325, 2.26387646045867,
  -4.63584947274609, -8.85519930079019, -3.74525746145642, 1.9813383447589, 
    4.60743921246128, 1.6105297186717, 0.173267125406393, -2.20588679277751, 
    1.28392207464239, 2.39675911670017, 6.46542418124481, -10.3161185510907, 
    1.18945056724182, 5.13960552857742, -5.7887274994311, -6.15174618988476, 
    6.11257068629742, 8.43772142844547, 9.76333403300334, 1.32488853223094, 
    -2.79190921460847, -12.3433019369319, -13.1082221517634, 
    -8.95483460679821, 1.04371691863926, 5.88891958523523, 7.08303382064151, 
    9.28595067859809, 4.230462578095, -0.914419784420183, 0.319074516238557, 
    1.73091692615695, 2.19219593171421, -1.13903590088191, -1.4200422667287, 
    -2.86096782449181, -3.54460608330933, -1.0802785459308, 2.93504584700959, 
    4.54149627870502, 0.816552927843327, -2.95255057735831, 
    -0.178751742737834, 4.20672377585403, 4.98744579605763, 5.770095048917, 
    0.687469529302349, -1.90215996153946, -11.4362793774947, 
    -8.62738809793247, 0.127891486256754, 8.79285751646247, 6.26370310615449, 
    -4.0524345050651, -7.54410467951377, -1.04387934339274, 
    0.970523580784417, 0.30043619051657, 8.46532917144086, 5.65961156535299,
  -7.00482564989271, -11.5109162566851, -3.05046997377207, 9.36667666073918, 
    2.43620464070772, 1.06145715277359, 3.1562652686034, -10.5453650063648, 
    -0.512033406384951, 2.31140255993605, -1.92177041949125, 
    -5.39888590224422, -2.36101565208505, 16.1414728989977, 7.02831108645299, 
    -16.4525893876982, -3.63850715950525, 2.72787822994119, 8.6060852713414, 
    4.09276005267346, -3.70479532702576, -3.49644378005062, 
    -5.74143911885609, -6.87154164786177, 1.22490657339169, 12.2696833231404, 
    6.58727111528933, 0.316013893611846, -3.926428080618, -10.7493144844848, 
    -4.08649690184961, 14.995101367908, 9.17160738005587, -10.2429690347904, 
    -2.72556646505816, 1.36652818730212, -9.29250596596726, -8.0296170471197, 
    1.10720668547312, 8.26303210418984, 7.32405165532348, -1.51728455474817, 
    -6.72694820516835, -3.60071813575427, 5.99472353737004, 10.9281667409664, 
    -7.06027355237811, -2.50886799204111, -1.11428767070458, 
    -11.3006983516569, -4.94544996289326, 8.34547460011028, 18.548586591372, 
    2.75232140505684, -15.7629887639928, -14.6715136378202, 
    -4.42781259923626, 3.91501205446889, 10.226983459724, 7.06257756488567,
  -6.83600810091251, -18.9386418037332, -0.66515149431171, 13.9526801947443, 
    -0.249177688361859, -0.262875518376207, -1.34501539948126, 
    -3.03102469681717, -1.23014198431497, -4.11635593295063, 
    -2.75549887669781, -3.5284507820381, 3.42043000153557, 13.2831466884076, 
    4.84934727743143, -9.05108413844223, -12.4413451544458, 
    -1.90384700311454, 7.92676080862972, 6.15264598392201, 
    -0.602309336049038, -3.04676350256767, -0.307403756370115, 
    -3.210715410992, 0.804213637980716, 13.6684483894639, 5.93627991272697, 
    -8.32944818432159, -8.42626995770758, -10.5180125953022, 
    -8.42017587919334, 12.606122687446, 4.23725452079239, -6.94335170813566, 
    0.851837224383171, 6.03289805414883, -7.1230927407628, -10.1927708170735, 
    3.22916331135034, 8.77009159798721, 6.37278854186292, -3.1766882962065, 
    -12.2419634825788, -8.45548097687739, 8.55608367579353, 8.2950195027505, 
    -10.2236092654721, -1.94680533822649, 8.46434072982048, 
    -5.83586787633268, -6.47933713659133, 9.19433922080085, 15.0078905127723, 
    -3.96712839634537, -12.8617980772345, -17.2369464262038, 
    -7.75570397767158, 7.62780115794763, 10.6967744450127, 7.19921522466462,
  -8.52584474614172, -13.6717467303138, 3.17528556770024, 10.1918425219369, 
    0.282913494064233, -0.930758822553884, -10.6530528336842, 
    -0.462440410164557, -0.729724098191994, -1.806704926941, 
    5.38764730997986, -0.0605376231137302, 2.01914990252989, 
    3.00228543971165, -0.50577454658424, -8.84848493098543, 
    -11.0242392545245, 3.75342972389416, 6.30174249767444, 7.30963611906546, 
    -0.500538843133897, -7.44390224978934, -4.23733790760242, 
    -4.43488136909298, 6.87023909221207, 9.68158593515028, 7.92464159735823, 
    -9.29354871159473, -14.4692235840524, -8.97726136527996, 
    -1.36899976051422, 4.73128190753313, 5.6227304043326, 4.44748054508678, 
    0.23604027020905, -3.74073240813528, -9.3246783793847, -3.43214994756306, 
    5.03804687012699, 5.60229706530684, 0.843673643487789, -6.56682420057852, 
    -10.4495406566888, -3.52489219981045, 6.83003632313563, 3.85461800270722, 
    -2.5833202494528, 2.23957919349959, 1.22565200995846, -7.47225572190618, 
    -0.183396179654662, 8.91164081310405, 8.23919897061974, 
    -2.42317947090945, -14.0462484265763, -12.5707481365768, 
    -3.74598262939814, 10.4356233295991, 9.09399092705146, -0.351424010133193,
  -8.28009034264433, -6.59336243342637, 4.30625504287454, 3.13691243538775, 
    -2.9720997812525, -0.174336677045915, -6.6860548272502, -6.633386913525, 
    7.9474124785795, 7.99170929420387, -0.0188217703028618, 
    -2.77977503566031, -2.55655834872181, -4.18907432508255, 
    -1.53781626369041, -7.12730123484396, 0.0655336267026161, 
    9.22626171140301, 4.5276225866491, 2.85908153889821, -9.45659942711179, 
    -8.14277847000871, -3.32818987732377, 5.09034459752886, 11.0428521582391, 
    6.47888598196899, 4.43456806287801, -7.06920473191928, -11.4644220083093, 
    -8.68253258721978, 1.45753711554549, 7.95424997502676, 9.71623682319055, 
    2.32168003212539, 0.107575383058157, -4.9575860443303, -8.64461291307045, 
    0.0700958747144502, 5.47110000102063, 5.88784215651554, 
    -2.73736858943605, -9.00210961461894, -7.68690725758101, 
    0.549068208897767, 7.37622805953734, 5.47683651356438, 0.755795985218712, 
    1.51738633049332, -5.36537346702348, -6.29036597774844, 6.23820557749546, 
    10.2955132214871, 4.42073153447871, -4.76483967056126, -10.3683723900419, 
    -8.06058779652053, 3.63342104854193, 8.48972289266175, 7.72164823675928, 
    -3.28444417881134,
  -1.53121523920967, -4.62021259171362, 2.78001080744063, 1.2040886586489, 
    -1.67940562998466, 0.475385800190039, -0.982001238209556, 
    -0.223610355184215, 4.39457402408205, 4.25444749932132, 
    -2.22475670124919, -3.40207604611028, -0.538587438072756, 
    -1.68924498440223, -2.26001405886649, 2.49055758049224, 7.23709420551312, 
    6.28320417057345, -0.472869319479991, -2.30534132151129, 
    1.07438656828001, -4.57819854769437, -0.645529588582966, 
    10.9495048705179, 8.13271225008029, 3.49979922512608, -2.8260036745703, 
    -7.49761696757705, 0.675810749562483, -0.91684467195347, 
    2.80502301041423, 5.46486550765168, 4.0104498792077, -1.48083998229161, 
    1.12915054782545, -1.74552674854567, -1.73853329439661, 
    0.859773732040356, 6.40492729096864, 3.40532684019005, -3.62515239647249, 
    -5.26746099558471, -0.786372466009375, 3.65349787023455, 
    3.65087696287946, 2.23805654611191, -0.0149159076563995, 
    1.54023618021769, -2.08778650518173, -0.893412790779656, 
    8.13207366803433, 6.49949472309789, -0.564627132262724, -6.0405137540156, 
    -3.01829517560295, -0.0410080647498436, 4.53268347725555, 
    6.79608897570458, 6.70923389968159, -6.75043787666718,
  3.57979151256103, -3.16299861184415, 2.64845456683819, 0.190246528604754, 
    0.548867280922564, -3.0724365400082, 1.89398326506956, 
    -0.502714493361086, 0.0611594697023056, 7.09093544665804, 
    -0.971161252920141, 0.616014838166878, -0.94634234753227, 
    0.253981004447517, -0.073420832294591, 1.63435049742376, 
    4.84591599821686, 7.25818333591938, -2.22775011346297, -2.44637809661107, 
    7.36004888502943, 4.7152013548772, 0.309813512693967, 4.74970812247156, 
    4.94438880528214, 3.45179575520717, 0.648506070008928, -4.17948279032095, 
    3.0092971647984, -0.684217063925533, 1.00836163506691, 4.20231982002294, 
    3.49573181071743, 0.758700197910439, 0.230377184425596, 
    -0.332262026727818, -2.09228536426974, 0.392096763363313, 
    4.33387590538393, -0.877085300990405, 0.096601124163225, 
    -1.27425955487862, -0.0527105194959604, 2.42999128407631, 
    2.55596707627893, 1.62944694562676, 0.139118672580841, 0.805341584591204, 
    0.131277189282439, -0.407658834616686, 4.90036329989631, 
    -0.164309792334153, 1.14905957339115, -0.85879654541533, 
    -1.08572860521934, 0.704014880629449, 3.72816123890704, 2.97226998736758, 
    1.11957463650563, -5.86061522086166,
  3.6947670463009, -0.090502644338625, 1.73805430681159, 0.703554800035053, 
    -3.2898834735668, 0.573424891245625, -1.92997351722276, 
    -2.81994391613589, -2.53600617799401, 2.05835233491843, 2.89243086178676, 
    3.51506669239874, 0.744329445313137, 2.29786342657671, 
    -0.218927281095255, 1.10933967096319, 4.99921974755525, 4.0090833794376, 
    -0.482271738681725, 4.33858347161848, 2.63379107557871, 
    -0.520745692095245, 1.90901723653691, 5.19002735717112, 4.44518019307144, 
    -4.40820384808655, -0.0197410193168409, -0.402118435390555, 
    -1.88861639495012, -1.37556539393769, -1.54829727284177, 
    -3.81694573628643, -3.56250189265565, 1.58581258703472, 
    0.153285220750812, -0.815326528825296, -1.03052649695663, 
    -0.112410063966847, 2.64919581058562, -1.1213448167276, 
    -0.425502750221477, -0.933356678879985, 1.78878790196917, 
    1.85320390218267, 1.99887458767234, 1.30470728176053, 3.2313888953044, 
    4.75997709400838, 2.64172341632193, 1.56288473098042, 5.18267393772354, 
    1.98542047366807, 1.19525303254459, -2.16474175177328, 0.148366952754004, 
    0.192205307731924, 0.165770891721897, -2.96882848375232, 
    -2.26141793962228, -3.55695359155954,
  -6.52745078974981, 2.98974459556686, 1.52182149632637, 0.674254417145973, 
    -2.07180180272488, -4.18670189276559, 0.885770748308184, 
    -0.0934176184585182, -3.81687820737151, -8.13757753308038, 
    -0.0253583233568414, 1.44610880373536, -0.534277065508913, 
    0.436839799669676, 2.93599217090046, 2.26116064647054, 0.369119028469098, 
    -0.14857280835952, -2.38452901992537, 0.635862408251428, 
    0.759316142182789, -2.37937889364785, 0.882785510666278, 
    -1.46054941072091, 5.0629216804441, -2.17768369394176, 0.128228854004955, 
    2.09092256456437, -0.980249784816398, -4.37029919198867, 
    -4.72425446354263, -1.82747645244111, 0.237688685087557, 
    0.0308995377523465, 0.40887111675468, 1.1305923940289, -1.5659072298917, 
    -1.47263588553979, 0.536099614888515, -3.79885464433871, 
    -1.51938442927571, -0.609967701521094, 1.35539407330033, 
    -2.5034484572096, -1.72695766878636, -1.48726815556102, 
    -1.66620691878808, 0.596817159944479, -0.442670304811151, 
    1.53921076491917, 2.59812564239859, -1.67476533302141, 
    -0.853534250451328, 0.0137418866363326, -0.209066066321769, 
    -3.39528560976309, -1.41649140078062, 4.97091085101864, 1.56964847843799, 
    -3.70340760811202,
  -6.5406206964961, 2.2147878826327, -0.39719068719951, -2.19125016297076, 
    1.4338767102325, 2.47976438987902, 2.08130109387511, -1.62329409206947, 
    -6.49723199395309, -7.08609632361568, 1.06067488544761, 3.15129490743564, 
    -3.00215902853908, -0.980733241833249, 0.133079040274066, 
    2.78919991180589, 0.768140274143033, -0.00360880849414652, 
    -2.96520676381572, 0.539715271568644, 0.0449888247704269, 
    -2.01792268386277, -1.42227008591771, -0.318479191781852, 
    3.31702255271546, 1.25931518040875, 1.42716725183521, 0.855971086635419, 
    0.899550586461357, 0.0539820565438335, -5.87108080931923, 
    -6.28411964494565, 3.15997122015789, -2.58849035351401, 
    0.390335607585448, 2.31398315215669, -1.49984844486215, 
    -3.02961418237044, -3.6359207242125, -4.21848569223975, -2.7419929932058, 
    0.990167916905565, 3.24909493438434, 0.556354197683402, 
    -0.685838621031647, -3.63930894734584, -3.17407303067404, 
    -1.24113946317876, 1.01073002439091, 1.13896273560604, 1.23751385919969, 
    -0.130036718070603, 0.0420962487853358, 0.600472755195386, 
    -0.243571334040344, -1.29245221577267, -3.91068490860718, 
    -2.98055057627079, 6.71870818548183, 9.08251374443724,
  0.565094833230726, -1.93217187707144, -8.14915084168082, -2.00742594671748, 
    4.5988770333888, 4.59689438435402, 5.36977110362504, -1.93323404823785, 
    -8.82829434181763, -11.9744514402183, -0.194729003807478, 
    8.04338941160431, -1.73482416570476, -3.00650245990687, 
    -0.463452861977118, 1.04651088117422, 0.459545326754207, 
    0.561313199776862, -2.70855279654968, 0.968289553601504, 
    4.16160202712056, -0.791289361119332, -5.6875606667703, 
    -1.71556266959999, 2.46897139452245, 3.58192258897782, 2.76886428057096, 
    2.33565045391606, 2.2919542649019, 1.64216222843091, -2.39097680569802, 
    -11.0502684530907, -2.06418768843978, -3.69138483543797, 
    4.72288857184472, 7.24447519518131, 0.903369102125769, -0.35993318589881, 
    -6.19738140326327, -6.84232562659482, -2.06179310897892, 
    1.98429054932759, 4.43166526770662, 1.60818477293312, 
    -0.0866698521811757, -1.58699817933862, -4.76127770973346, 
    -3.52824770885495, 1.63730482477438, 0.180662508468975, 1.06675942319265, 
    1.95332448438566, 0.646564518312003, 2.50970943095237, 1.96046253886267, 
    -3.093564940932, -8.34985239634545, -6.67869883624808, 7.52543057986676, 
    9.06167711657639,
  13.6582791264747, 2.47846757434715, -10.3619383577481, -9.42648721789218, 
    4.30047002334107, 11.5238992813215, 10.4510414096031, 2.03009847537058, 
    -6.53727967049383, -15.4861789832886, -9.44428952346337, 
    7.50474752069414, 6.94757172657607, 7.10315156549507, -0.260205486728304, 
    -4.92168043349928, -7.03758499948351, -1.04746686508362, 0.8419790399802, 
    5.89729135069114, 5.817537723839, -1.38550399386213, -7.96265535972788, 
    -3.75817520130749, 3.3644379534061, -1.88241735079166, -1.86792594514672, 
    0.497812287330304, 6.94422007079328, 6.05418597160593, 3.74715867601901, 
    -6.79286805548902, -9.20928064744118, -4.16303557023292, 
    4.96007188715275, 6.37308886470308, 0.919570935718915, 3.02991222524231, 
    1.03488199907009, -4.34397158062007, -3.09563587676096, 
    -1.71549689074449, 2.90816150397514, 3.79320558903042, 0.710004414039221, 
    4.53661904234701, 0.3901366188747, -5.66323318662082, 2.23759572438597, 
    2.7095625856579, -4.32694662503798, -3.93817832440274, 0.601606687806136, 
    2.02944691862029, 2.85078116706516, 1.63266365269916, -5.97957640501947, 
    -7.55616121768989, 1.61276797480961, 7.81509511678344,
  16.0992404467035, 2.76732755002009, -2.56433438566862, -9.77816100517961, 
    -0.253216616891402, 13.3901051141657, 5.56825332167319, 1.32034747641075, 
    -1.89676677605719, -10.9307883285183, -14.2080809451068, 
    3.10515510301705, 17.8683156309499, 16.2612704336111, 2.6660318707958, 
    -9.18239819209088, -9.54020909612614, -1.8857578781462, 5.85848314382934, 
    9.10210384414468, 9.52017937901306, 0.410994495061781, -12.2188240536066, 
    -9.89333590220254, 4.46154602005486, -0.248482297021874, 
    -5.9774280016471, -7.30066116252953, 5.90940819864558, 9.23693632724976, 
    4.96104143566737, -0.155151286216017, -6.77199266933137, 
    -5.63093627073198, -0.749559112858359, 1.24391182261474, 
    6.21484427628851, 4.70751357904153, -2.36584112924838, -2.05841211921094, 
    -0.161405326453607, -2.97123089119981, -1.87973181463237, 
    6.17524888940393, 3.4414954605437, 0.140952955615272, 3.4596118551708, 
    1.54077158291757, 2.50345669740604, 7.0558915193233, -1.8218789424532, 
    -13.3868947873869, -5.37760310549013, 2.14954782955262, 
    -1.57537455678595, 2.0150775225794, -6.53859095630163, -11.6724618035603, 
    -1.60696045332983, 15.2091704970771,
  6.03800188900061, -4.14729089067785, -1.87025829775354, 0.043780021075651, 
    -0.418671351692227, 1.55365622993503, 5.27458686889482, 5.39175230032009, 
    -1.84729873732889, -10.9347927382529, -11.1828851064118, 
    2.78487804379494, 16.9019638910521, 15.6404898467914, 7.06495669201165, 
    -9.45285978878509, -13.1763791710324, -4.76103864534826, 
    8.94325399094061, 13.6083493198599, 12.1529307421397, 4.46969923829883, 
    -9.80811802125958, -13.7174538756777, -2.43961613048613, 
    6.44526903082149, -4.46506808830363, -5.0143330664678, 6.34896719143943, 
    2.12606071611487, -0.376176087000431, -0.929063682323387, 
    -4.04745765357732, -5.78567344395998, 0.908212894497921, 7.7775843720504, 
    14.1848741489685, 5.43193539790937, -8.42053688521199, -4.19509081172413, 
    2.54881038480405, -4.1060138289057, -1.24027423724495, 6.06046004091299, 
    7.65150733080205, -0.745836964629857, 0.984499956885733, 
    4.09388267867798, -1.16343633635427, 2.80887563857139, 1.70301791012592, 
    -12.4441861645017, 1.47083795908898, 3.35257555891404, -9.72277714276913, 
    8.70941588432953, -1.84330430584944, -9.72880248900151, 
    -6.82943715783329, 10.5619308693579,
  -9.08890593333562, -6.01777997480791, -3.56399933356887, 1.38829775530378, 
    4.60265028400796, 5.19343515477939, 12.7942942913669, 3.88715906067078, 
    -6.79163419248196, -10.4053540507782, -6.76051156346249, 
    6.66260951572253, 9.23830029683243, 9.61181447337688, 9.75496626856395, 
    -1.04327557049881, -14.1748052866045, -10.9183746110816, 
    2.60775363938876, 9.65967307148143, 10.2144637887382, 2.68615012541231, 
    -12.2630468813757, -11.6270157182227, 2.30165107139568, 8.36079182916909, 
    1.08026305836567, 6.7312215274332, 2.56992095169326, -3.79788631607596, 
    -5.44797863537115, -6.57186332969127, -4.54071571597575, 
    -3.11137503826381, 6.13944577181252, 10.4758583596871, 8.64362027744198, 
    2.00381140193089, -4.07340765643994, -5.89726247691269, 
    -1.26460229437324, -10.1932229866945, -0.699825882552561, 
    10.6944466534455, 13.423221144035, 3.5882712885991, -1.02891585653616, 
    -5.90376049360133, -8.61717323573547, -2.93103814810464, 
    0.0943383736634004, -5.35041492308317, 6.89009152234918, 
    4.92673597719531, 3.01652792563349, 13.8321032246128, 2.40152683019023, 
    -2.66317117339772, -8.84702929026601, -5.02485206979732,
  -10.4049123955188, -4.74991764544967, -0.372390790695416, 
    -0.241270563917005, 5.62540170016186, 8.12516650615211, 4.29591641140499, 
    -4.6168019317038, -4.94113912272139, -2.8137497441032, -1.03203762570508, 
    6.54556595591892, 6.3399377366424, 5.49949576720346, 6.29030189850766, 
    -0.8627484278553, -8.19154007505794, -7.79487190706501, 
    -4.77630792265743, -0.489378775032945, 0.22471615397676, 
    -2.56613973703453, -8.54809806238157, -2.77564134084454, 
    8.37375860771824, 5.67601340638984, 8.02674165583649, 9.14754591203777, 
    -1.82534637583664, -0.719564512117791, -4.39598582564017, 
    -6.11841006756343, -2.44005949454842, 0.900308137217475, 
    5.52169705866377, 4.44833986685104, 0.0308849639261374, 
    -5.23436792546687, -4.69323886955685, -8.03786767071338, 
    -7.36920116014356, -3.78160334492942, 4.09000137506903, 15.1613175989845, 
    10.6880087241307, -0.404667734587072, -9.81985886808948, 
    -16.5297055988129, -6.21073905109818, 2.6797784278022, -3.48390584155067, 
    -2.54094961947363, 3.42290110388965, 7.88918598029895, 14.2558422727073, 
    8.95987914193951, 4.19960010692016, -0.923677597321415, 
    -7.62779556359521, -8.70433062275619,
  0.568511501269831, 0.281738613467411, 0.92177104680294, 1.27532671805745, 
    2.78516709697503, -1.42829435434583, -6.44595993642938, 
    -5.47440306205589, 0.606505802174156, 4.09769177005636, 2.79091350789308, 
    4.72594074679191, 3.5140464770363, 1.36368531982318, -1.05560213979481, 
    -7.50491351951956, -6.3443234793713, -2.31561217056731, -4.2822074283174, 
    -4.39169073003945, -2.01295125918763, -0.490718634110127, 
    4.40187951594881, 3.81408093135829, 3.74962268955555, 4.52738199362324, 
    6.90900012576798, 2.44588555986686, -0.530455811300957, 
    0.456625450785844, 0.677672460578931, 1.2380483181918, 1.82545142754429, 
    1.60289660689775, 1.85283553951963, -1.32281232762078, -8.33021313741466, 
    -13.2255937293582, -5.87444448356849, -3.55739027959986, 
    -4.42010671561636, 10.9461227455091, 11.5882029689301, 7.80265846938543, 
    1.42908248833993, -4.58605415005487, -13.929470044171, -8.24695496082125, 
    1.14939747802777, 1.30578656465706, -4.91237954284266, 
    -0.635508576867734, 1.99504263123834, 4.60599054762536, 7.21889402980788, 
    3.99763437282036, 6.70409443169112, 0.219433244818976, -8.71571205321212, 
    -8.1776360996,
  3.01749942948141, 4.68240391488321, 4.47467428649546, 5.3071291479493, 
    1.82505744263389, -4.12206366818579, -8.90017567994595, 
    -8.13463321941018, 0.131135364292304, 5.43694774014763, 3.91944187342193, 
    3.61831898481206, 3.10910935542225, -0.618478882099131, -5.6674465747795, 
    -9.79708911429074, -8.08602762522344, -2.48938039028236, 
    -1.19318838873002, 0.00694448142492064, 4.55779573378088, 
    5.78663979588877, 5.64358577496637, 4.42294834131557, 3.20395338367797, 
    2.57738747183791, -0.0637039516452208, -2.55739339941335, 
    -2.47918154009513, -0.824361011535635, 1.47765818312938, 
    2.46991696627624, 1.47252777174753, 0.168231975630355, 2.04744742013706, 
    1.24773131811952, -11.7358966402817, -17.9016930046314, -3.9768672496424, 
    6.00962614625325, 8.74930437249402, 14.9585230954767, 9.7823545319751, 
    0.659613350096675, -1.50126459611281, -6.10478587555804, 
    -9.21968520673323, -0.778561988479015, 3.88072934674314, 
    -0.0350861019728684, -1.2734707158754, -2.81846888496291, 
    -3.6156545536635, -0.129702406308316, 1.89997988374196, 
    0.750969221017815, 2.49128061489011, 0.559538968226209, 
    -6.39057630343191, -4.88379789508208,
  0.0373437689152269, 4.21892054963698, 6.38498335465194, 6.73771054240844, 
    5.31638982113985, 0.838008414156993, -5.59140325323673, 
    -8.84611321051935, -6.17919474138623, -1.20477789180962, 
    1.80756981642166, 3.37755399319123, 4.031813941612, 1.1347458969967, 
    -5.30377643919804, -9.75762851234351, -8.15654132671122, 
    -2.8912245030581, 1.99271081359576, 5.05026675857359, 6.33225347070439, 
    6.38470703862092, 6.05260781479026, 5.50337724929123, 3.81799098503674, 
    0.785384814402459, -2.38192287311423, -4.51736827633253, 
    -5.07338883007623, -3.39260219570392, -0.601796242098797, 
    -0.544756367046579, -3.53828789761248, -2.75848365092672, 
    4.57402223138865, 7.59014155724339, -2.50008405113121, -13.7502123932993, 
    -10.2052860429622, 3.2994473532737, 11.6686870087359, 12.0080069977267, 
    7.80624619712314, 2.02113749548186, -2.39557493610879, -4.12029471268078, 
    -3.73438214793995, -1.21525137823036, 2.9884612925858, 4.27029857197315, 
    0.631419904648731, -2.88964503616766, -2.21903692303056, 
    0.24500457046989, 0.722527100124814, -0.64240710253231, 
    -2.14762192391768, -3.59146265847274, -4.66226399535471, -3.72436100698875,
  -2.63638327896604, 0.235273397428973, 2.75558907834126, 4.83338847556666, 
    6.13259997028203, 5.61666271544753, 2.38175817863231, -2.76161350069635, 
    -7.03488536752258, -7.81390454345622, -4.98578229863087, 
    -0.900339782683934, 1.78107149807855, 1.74125494028777, 
    -0.524934420638794, -3.21735979092572, -4.20806028365935, 
    -2.43154703703225, 0.945764061630278, 3.77621823094461, 5.05889050122699, 
    5.26756564266923, 5.23288606299506, 4.84807861890975, 3.17746019307084, 
    -0.160365476187043, -3.9764829985377, -6.08336968989958, 
    -5.20690788959916, -2.56539987469275, -0.865665593519049, 
    -1.32372919638903, -2.09368729065129, -0.263171730212354, 
    4.27310586984676, 7.56692102357522, 5.47803078866303, -1.35287682386763, 
    -7.18884934051504, -6.53011102924768, -0.8968766743017, 3.53732303332624, 
    3.50824189302733, 0.656692050861484, -1.59589055632941, 
    -1.44670156046803, 0.465145222704983, 2.14809584270656, 2.21280261822334, 
    1.43368515831616, 1.24604077288933, 1.84914035420667, 2.69911025776139, 
    3.24583050996973, 2.8838678123262, 1.08576107397962, -1.95997512202037, 
    -4.96772068583549, -6.26322644111405, -5.20360503852571,
  -1.64879007409176, -0.798613923001449, 0.793284366838634, 2.55315619214473, 
    3.71432896813913, 3.60585943761591, 2.04296297171458, -0.55983086147991, 
    -3.37034917045459, -5.39499514252008, -5.84863678409686, 
    -4.58603332948039, -2.29826987350408, -0.112675488948251, 
    1.02209974958183, 0.780268849435938, -0.418317276077301, 
    -1.62744439157869, -1.90578769542616, -0.979607818584794, 
    0.622564529967407, 2.04205214333873, 2.60114648454128, 2.1241389786587, 
    0.961271823313385, -0.243831474242633, -0.908903307712667, 
    -0.868619269977864, -0.330169029658417, 0.410813611282111, 
    1.10981552373522, 1.63461086628442, 1.97812166228208, 2.18755707520817, 
    2.28613763505671, 2.15084089231284, 1.55262776900878, 0.403892975311253, 
    -1.15409004384029, -2.8492010871959, -4.05196514466307, 
    -4.12923874805799, -3.11115139571384, -1.63766781955518, 
    -0.453248556948902, 0.0193505337845474, -0.156949777726865, 
    -0.543087033930112, -0.636006031067208, -0.180726114888346, 
    0.774064915743921, 1.99705302134099, 3.08308995844681, 3.6845733532883, 
    3.65518192147301, 3.01519780461155, 1.92195203438333, 0.611997552506368, 
    -0.659012870246424, -1.54491756339169,
  3.57809814137005, 2.73016887481485, 1.69923011063025, 0.615201558693873, 
    -0.405882227968683, -1.26750608002501, -1.91245471757324, 
    -2.31144515292934, -2.46386749059022, -2.43407850851568, 
    -2.31965721893497, -2.19754513477629, -2.10195532178838, 
    -2.05053568761681, -2.05170518555856, -2.10025663331724, 
    -2.17122194417088, -2.21768917302806, -2.17390142812651, 
    -1.96122973861701, -1.50607101111061, -0.780826998507698, 
    0.1848107982262, 1.30720223534257, 2.44522158135528, 3.42827836246349, 
    4.11256476114653, 4.41693339622388, 4.30593575397504, 3.79259749657995, 
    2.94726995318406, 1.89049378392714, 0.763814846663309, 
    -0.300190263882543, -1.19496132936246, -1.84404333080437, 
    -2.21956264197925, -2.33427407027989, -2.22280455245184, 
    -1.95436278965718, -1.63874956161866, -1.37835056204587, 
    -1.22459375092764, -1.18118661404781, -1.23481208934715, 
    -1.35676055537885, -1.49509908689718, -1.58291437532138, 
    -1.56453092237116, -1.3868846890696, -1.00832036299097, 
    -0.430600538766631, 0.337797095926045, 1.24366296047621, 
    2.17933456459081, 3.03028066818582, 3.70904631696222, 4.15541665370669, 
    4.31393748955354, 4.12696329872311 ;

 time = 14.5 ;

}

