netcdf filter_input {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 10 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double concentration(time, member, location) ;
		concentration:long_name = "tracer concentration" ;
		concentration:units = "mass" ;

	double mean_source(time, member, location) ;
		mean_source:long_name = "mean source" ;
		mean_source:units = "mass/timestep" ;

	double source(time, member, location) ;
		source:long_name = "source" ;
		source:units = "mass/timestep" ;

	double source_phase(time, member, location) ;
		source_phase:long_name = "source phase" ;
		source_phase:units = "radians" ;

	double wind(time, member, location) ;
		wind:long_name = "wind" ;
		wind:units = "gridpoints/timestep" ;

	double concentration_priorinf_mean(time, location) ;
		concentration_priorinf_mean:long_name = "prior inflation value for concentration" ;

	double mean_source_priorinf_mean(time, location) ;
		mean_source_priorinf_mean:long_name = "prior inflation value for mean source" ;

	double source_phase_priorinf_mean(time, location) ;
		source_phase_priorinf_mean:long_name = "prior inflation value for source phase" ;

	double source_priorinf_mean(time, location) ;
		source_priorinf_mean:long_name = "prior inflation value for source" ;

	double wind_priorinf_mean(time, location) ;
		wind_priorinf_mean:long_name = "prior inflation value for wind" ;

	double concentration_priorinf_sd(time, location) ;
		concentration_priorinf_sd:long_name = "prior inflation standard deviation for concentration" ;

	double mean_source_priorinf_sd(time, location) ;
		mean_source_priorinf_sd:long_name = "prior inflation standard deviation for mean source" ;

	double source_phase_priorinf_sd(time, location) ;
		source_phase_priorinf_sd:long_name = "prior inflation standard deviation for source phase" ;

	double source_priorinf_sd(time, location) ;
		source_priorinf_sd:long_name = "prior inflation standard deviation for source" ;

	double wind_priorinf_sd(time, location) ;
		wind_priorinf_sd:long_name = "prior inflation standard deviation for wind" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;
		location:axis = "X" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
                time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		time:units = "days since 0000-01-01 00:00:00" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "no calendar" ;
                advance_to_time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		advance_to_time:units = "days since 0000-01-01 00:00:00" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
		:description = "Saw tooth pattern for mean source at grid points 1 3 and 5" ;
		:model = "simple_advection" ;
		:destruction_rate = 5.555556e-05 ;
		:history = "same values as in filter_ics r3002 (circa July 2007)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 concentration =
  4924.10747884102, 4172.44107017966, 3405.82353170351, 2838.91189156883, 
    2574.63559485657, 2299.77454361968, 2026.6312412118, 1886.07056314528, 
    1764.6490788102, 1657.27114789251,
  4945.69096625066, 4173.23666925717, 3328.71554246707, 2846.17239358214, 
    2577.60084708482, 2275.73235173497, 2070.33108080167, 1917.67032530519, 
    1771.29497467247, 1690.75025584681,
  5018.88972761714, 4106.6014394109, 3412.84290410569, 2906.52180390099, 
    2505.83916340037, 2254.77391565149, 2041.58593644403, 1937.34658857106, 
    1781.26595310229, 1666.8303314331,
  4966.57751625612, 4116.5783512006, 3352.63672107293, 2886.01603089924, 
    2566.01282428024, 2254.23359284475, 2065.9244308836, 1899.92336820227, 
    1775.72145118492, 1655.47171264901,
  4894.80361667694, 4132.28353488566, 3335.50535553369, 2898.90465201079, 
    2532.17470018573, 2264.86799764488, 2060.31909636037, 1900.50829531702, 
    1740.13270431707, 1661.26867837486,
  5028.6694330573, 4092.11358538244, 3383.50724828674, 2838.66284803882, 
    2532.98054008453, 2225.59985719235, 2021.6671653032, 1913.14589339301, 
    1735.89053054651, 1652.99225235236,
  4925.51290327203, 4103.06829804821, 3431.76318221917, 2924.39176545205, 
    2534.04516633297, 2260.9501391778, 2071.56434890848, 1944.22839067543, 
    1757.38801529808, 1662.33300326783,
  4983.01239556323, 4133.0382043153, 3373.208964453, 2876.82500831065, 
    2592.53924495123, 2235.21053006339, 2027.79402812407, 1894.97913895726, 
    1778.82909894927, 1652.26922646599,
  4915.97324539543, 4180.24894646556, 3367.37972692498, 2841.92042918964, 
    2561.33526062596, 2269.16533837797, 2065.32104356297, 1907.29727737165, 
    1778.36888243111, 1668.63328179326,
  4931.09176697597, 4190.08773460702, 3342.27474504449, 2921.49147295283, 
    2576.38719554849, 2261.94387954176, 2039.90458302071, 1915.91243317584, 
    1778.22938018388, 1667.91096949921,
  5019.78917516078, 4085.97217592396, 3375.51687689946, 2868.31907130621, 
    2573.48115301356, 2264.42756643888, 2051.5373398129, 1915.49504971136, 
    1773.34882732472, 1675.59389507398,
  4924.36612456836, 4126.07629097544, 3390.26448218447, 2911.6426612775, 
    2557.2799787717, 2223.01223380153, 2068.68384854592, 1909.50110377618, 
    1770.4178894942, 1673.55602278965,
  4859.71220814277, 4121.18746414821, 3318.63056508771, 2843.02357158759, 
    2552.48835019096, 2304.02613525355, 2044.91962874357, 1909.28034923807, 
    1767.06004670869, 1654.92069355955,
  4936.59518068566, 4125.75160696811, 3377.16073304764, 2839.22921620396, 
    2583.27420112754, 2276.94178514069, 2042.02212782508, 1903.04652128871, 
    1752.72107001841, 1674.09417676217,
  5104.66650349754, 4138.58355386587, 3392.9602576871, 2899.49859656006, 
    2557.97066793503, 2224.16594828241, 2040.61019627005, 1913.78765964501, 
    1783.83726968603, 1663.95924742126,
  4891.4506511284, 4116.08348629678, 3401.79021858421, 2900.42981268785, 
    2564.54295074198, 2242.42225672859, 2052.10150889734, 1908.51309281453, 
    1765.12663479853, 1679.99144486292,
  4996.69557948961, 4147.40958095827, 3347.65527699646, 2933.34895679199, 
    2561.10465702598, 2287.61536415957, 2063.66764406863, 1893.06316643151, 
    1761.60743117224, 1660.60173243095,
  4978.04851021947, 4132.19940484389, 3328.1223336241, 2851.31589754639, 
    2625.69370318132, 2249.61771428419, 2047.44154538806, 1890.81050942142, 
    1763.95042456331, 1667.22189752151,
  4902.61374855636, 4163.4330130031, 3393.70609611685, 2843.04095838105, 
    2536.62945452891, 2231.90100654581, 2058.15387141905, 1908.46252313845, 
    1763.08379726238, 1670.53269037302,
  4975.85787254064, 4153.90000476752, 3345.53877783797, 2951.14268211444, 
    2518.20062893968, 2277.33619439965, 2068.81244966285, 1883.0612854159, 
    1741.26003780002, 1662.0554482122,
  4925.56148826297, 4121.97174580343, 3355.2089565169, 2829.78157831064, 
    2515.43416787498, 2243.89498497764, 2033.71640577626, 1913.52517373455, 
    1783.58259578713, 1683.89928795636,
  4853.63846890152, 4119.63534417543, 3404.0387177831, 2948.7277477238, 
    2573.54010094723, 2242.67005926766, 2062.17965324251, 1895.04340887177, 
    1761.58071547995, 1660.26324201232,
  4937.42824047194, 4114.91200627061, 3331.07837525047, 2850.73195893742, 
    2572.60333887499, 2249.67828643074, 2058.22458193245, 1934.859843034, 
    1780.39782019586, 1663.36077067953,
  4992.48944463925, 4118.79305180575, 3384.5042757799, 2869.59950287399, 
    2568.18779953661, 2258.91826580279, 2119.86962119204, 1898.36482943309, 
    1757.02915846728, 1665.88405735656,
  4975.29337339233, 4123.77377180451, 3338.26576372866, 2915.61898402916, 
    2505.5834679552, 2261.57544374214, 2057.82117699314, 1901.05054811384, 
    1780.32714262305, 1665.94971084014,
  4907.16056447814, 4110.36297796599, 3401.13569543261, 2858.85899986819, 
    2580.79615970831, 2294.62174228986, 2053.58934029893, 1894.79280058124, 
    1748.69413753122, 1676.10335460623,
  5017.01561239787, 4128.24168454176, 3375.73967887497, 2899.18878728708, 
    2557.42248741468, 2290.48449420282, 2085.40656178656, 1907.97603516998, 
    1757.74085999859, 1660.390888009,
  4952.91974591395, 4118.7094496836, 3350.40797717644, 2918.79316919046, 
    2575.72634722533, 2246.81201977311, 2039.51270815812, 1904.99517229271, 
    1765.8265989734, 1677.95221387727,
  4958.47183276314, 4105.29944764028, 3390.94430977458, 2880.221587193, 
    2576.33683577496, 2277.09242027693, 2063.86521766816, 1894.11844338017, 
    1757.6818355244, 1677.62818213841,
  5011.95929963519, 4105.46479102706, 3386.14557420067, 2875.78126097136, 
    2556.62437554087, 2248.25501831408, 2058.77117082383, 1886.44684752908, 
    1752.43276982282, 1664.2567686023,
  4941.21271360704, 4145.52685300221, 3330.1601323144, 2912.33678416362, 
    2520.81219995364, 2269.92292177755, 2046.59018431679, 1902.30096124077, 
    1794.61455500601, 1657.61638212371,
  4938.81803859002, 4112.02860706954, 3377.21251033578, 2856.67324882303, 
    2619.63666097746, 2250.54111352806, 2018.73942091893, 1906.56028787748, 
    1765.78826800501, 1662.39787960053,
  4899.09933467281, 4161.17464263595, 3341.84348274926, 2854.59683873369, 
    2565.4147075227, 2253.32873358592, 2060.2337022076, 1874.91431591569, 
    1774.76384443292, 1664.98683767947,
  4980.36985221169, 4121.419368115, 3389.46092056523, 2885.1716603269, 
    2551.66979999718, 2276.01185732799, 2058.83043949485, 1885.00103991941, 
    1768.64837676502, 1671.22387771715,
  4943.48753676914, 4121.83380769119, 3381.10284955992, 2845.68624026062, 
    2560.62572655083, 2290.4150001299, 2051.62188533585, 1929.04788744435, 
    1774.19371568002, 1678.63078111753,
  5028.7691412915, 4150.75652005708, 3361.63287047426, 2882.87003541535, 
    2593.30105435639, 2282.3994080671, 2068.66455244974, 1915.29894353838, 
    1753.22288882955, 1646.43793827731,
  4922.46419411394, 4133.17352322015, 3385.34390896628, 2892.28348232654, 
    2556.45990644102, 2274.62798221341, 2058.88829145113, 1897.82345072168, 
    1750.93477675961, 1656.04628028212,
  5010.43566262945, 4196.68826117273, 3342.14004290726, 2886.93709160578, 
    2554.77770211021, 2270.25596723217, 2065.7658697244, 1910.51792770547, 
    1753.20645706102, 1662.00586494342,
  4950.66002398226, 4133.39591317974, 3347.29950312946, 2873.1009747621, 
    2593.68005402925, 2263.7882118178, 2067.52310530651, 1884.80788613915, 
    1797.86127664701, 1678.02778967949,
  5031.67991513547, 4107.11549875191, 3364.56831812143, 2836.78139924309, 
    2573.16972360593, 2254.76268290576, 2066.05345563047, 1900.59224830643, 
    1751.00325150334, 1654.02334871879,
  4923.47087737786, 4073.68238368775, 3340.32276085659, 2854.21783112149, 
    2577.21352210948, 2265.89461673654, 2045.26989281491, 1939.92050843345, 
    1757.76358135731, 1661.3531148252,
  4884.34655116996, 4148.46450596102, 3310.08738996756, 2884.12254518231, 
    2522.26109594398, 2276.66604214414, 2059.09303695301, 1916.65065335011, 
    1741.04826881118, 1664.50008456896,
  4869.35421913921, 4135.42062500852, 3369.70381717181, 2920.5348542249, 
    2584.39594198427, 2247.5940401965, 2074.88991041728, 1921.21280592651, 
    1770.86300818709, 1673.27148681218,
  4994.68908470346, 4085.54067372871, 3339.41050631466, 2860.09202505971, 
    2595.50550551398, 2253.27809797025, 2031.62241488071, 1908.18992345145, 
    1767.07159542445, 1675.86607126328,
  4899.14833338372, 4191.66775299227, 3381.3417073612, 2877.531153253, 
    2542.07948231479, 2283.13425410869, 2034.4647376483, 1923.79068774272, 
    1769.55672485894, 1665.70507352318,
  4998.59023773509, 4102.3142366955, 3364.49411712261, 2868.39297949002, 
    2530.24102375752, 2234.66141885264, 2075.95192253843, 1917.7246371189, 
    1758.44293791255, 1663.68215839921,
  4919.61801633613, 4170.48034209738, 3338.71072040714, 2914.18316553297, 
    2583.41214167672, 2276.79697967736, 2057.45775150472, 1943.71071830189, 
    1779.42206689342, 1677.32081485733,
  4885.15551120383, 4221.15004185245, 3418.57942419492, 2860.24671540387, 
    2581.90729003953, 2270.46894912971, 2038.30273376415, 1903.97473672012, 
    1760.23464418901, 1653.25303990837,
  4956.80430752871, 4173.42894097739, 3327.38761219303, 2856.29906558697, 
    2578.13661884669, 2263.23592443515, 2046.89864519254, 1896.44419648505, 
    1767.43524267692, 1663.62445608896,
  4993.01946346254, 4124.82298167553, 3399.81848221031, 2871.47378438803, 
    2545.72608509745, 2310.19660258556, 2057.82415998198, 1897.75317673644, 
    1762.98273656249, 1675.34899444374,
  4943.45832922369, 4151.7435465293, 3331.47937582467, 2932.54404529082, 
    2583.34877989132, 2267.1426818812, 2027.93976711407, 1921.67116874386, 
    1767.29401929997, 1671.04639959385,
  4889.72596752956, 4161.83392757093, 3325.69927214453, 2905.13815582183, 
    2561.50632734598, 2273.25971814589, 2066.76374494633, 1914.7745659772, 
    1768.06602737415, 1662.73497886399,
  4952.58435892724, 4145.55735170017, 3364.50359743248, 2895.61720020222, 
    2544.33504028843, 2238.85469890697, 2034.83335547715, 1922.62627332099, 
    1754.02124586639, 1648.82040436274,
  4962.17043390543, 4148.58775588593, 3403.65935455951, 2870.40733480894, 
    2561.76085438, 2291.89904994417, 2035.38076671815, 1901.70035385103, 
    1760.05837529015, 1677.92464596791,
  4917.89486224179, 4152.15648266556, 3392.96106299889, 2845.78517452297, 
    2530.93726285211, 2234.66236560047, 2027.7236351859, 1871.56660475831, 
    1742.28058554082, 1669.55142383126,
  4907.13513833003, 4172.59098051484, 3368.46212837349, 2858.89761837634, 
    2536.54128908479, 2239.55665925984, 2077.9188651432, 1902.54358240741, 
    1772.54843969238, 1672.43677579623,
  4962.06623699868, 4138.68423860068, 3360.05339104016, 2878.97283131822, 
    2550.81626726974, 2232.76032162559, 2053.40256584139, 1915.99185414082, 
    1774.10634733503, 1661.59617669548,
  4893.02504977553, 4171.67245716942, 3421.94845442863, 2886.54116342041, 
    2557.16128097573, 2254.76836932528, 2070.65164938321, 1912.17919078047, 
    1776.06704219376, 1682.72606989297,
  4880.70535687378, 4155.49433753286, 3377.62302377112, 2903.68892981062, 
    2586.43029159355, 2240.10558871762, 2021.99981449493, 1898.4067403842, 
    1760.4087985369, 1677.02788748293,
  4988.09915220578, 4098.81798566761, 3357.91260397772, 2881.48514274626, 
    2520.80002825177, 2231.59256436541, 2037.09234296041, 1892.28930082294, 
    1763.74837332099, 1670.67462478152,
  4973.05408692204, 4168.76513668707, 3351.7854068872, 2867.86004334045, 
    2527.25133582989, 2262.59866471665, 2042.20277261294, 1913.78439773544, 
    1778.17461115178, 1668.73449136595,
  5012.14261512954, 4130.77364082642, 3366.49271760605, 2910.23678338535, 
    2596.15035591918, 2269.63364378325, 2048.0862392949, 1889.09558853009, 
    1770.2436377861, 1685.5429399133,
  4955.69153751345, 4138.02850020382, 3381.29595612669, 2853.01257245954, 
    2552.50982682736, 2234.26751802829, 2062.66599190253, 1959.96217312476, 
    1738.3342445704, 1659.42914913393,
  4935.64972334653, 4198.74670674874, 3331.0243468263, 2897.71441763406, 
    2574.13836579688, 2244.82822085188, 2057.00477997307, 1922.59890133151, 
    1787.03576821983, 1654.39880673335,
  4925.20486027858, 4124.75532094236, 3415.89507463518, 2837.52496374413, 
    2569.87792687266, 2268.63911222659, 2090.40229436239, 1902.60455960025, 
    1774.33025197419, 1670.08948463948,
  4947.98249414298, 4132.44157254503, 3404.87798385271, 2859.77667652408, 
    2558.9215812267, 2251.4354386069, 2076.84335399465, 1921.17195964298, 
    1763.13963572921, 1663.82500968443,
  4912.97773156659, 4157.64708360388, 3359.73610025199, 2853.69654919547, 
    2543.87892647122, 2253.37468820243, 2089.75988163569, 1902.65136632934, 
    1788.49243693174, 1677.82831313483,
  4960.26929934352, 4099.52800191491, 3368.39053365179, 2873.72056309179, 
    2608.05770335496, 2283.22580031984, 2041.86650668811, 1895.70713402126, 
    1752.42445678911, 1658.95033792214,
  4963.84449222548, 4086.48198096602, 3356.07002446581, 2900.40571718004, 
    2532.86026521758, 2256.75036406472, 2049.91945458839, 1901.6545473668, 
    1776.07781223255, 1674.90998026447,
  4985.45621860065, 4050.17748307422, 3346.722877817, 2875.99947957241, 
    2555.67344537599, 2216.38103501076, 2061.90046862793, 1900.05777197548, 
    1788.36475104317, 1681.26388684291,
  4945.74270050327, 4166.19837743956, 3348.00705478628, 2923.99931564633, 
    2603.82239229326, 2226.69431208587, 2055.26038532474, 1891.68720988837, 
    1753.2041817695, 1658.92143782824,
  5002.65039375406, 4150.92113117939, 3387.99274025257, 2862.10366385295, 
    2578.73711141712, 2267.44580470047, 2101.44867390363, 1936.67261530694, 
    1781.68133610382, 1671.14024211009,
  5001.20548716547, 4087.24184831794, 3320.4441439802, 2882.36415829933, 
    2533.82988755219, 2290.67053108295, 2051.83405874161, 1874.83865039907, 
    1751.16396888718, 1661.07758246947,
  4953.07708030152, 4154.56647076379, 3329.67514117504, 2875.60885348524, 
    2576.47905564425, 2224.52008060599, 2073.46531142399, 1909.48484908233, 
    1741.23174613839, 1659.48254464893,
  4961.21452977031, 4152.54088223782, 3355.08811550942, 2874.24031929228, 
    2558.08313595695, 2232.96058903707, 2041.50746537555, 1900.34536828054, 
    1757.50499681032, 1656.75821561953,
  4973.46925342563, 4134.44191159373, 3359.8922694744, 2858.19337681848, 
    2560.57101584645, 2256.0206193408, 2034.35422144698, 1887.09009069168, 
    1753.01973488181, 1673.06183834554,
  4919.18892047265, 4147.33044075448, 3359.83241187469, 2894.59213458651, 
    2563.30670668979, 2260.20636485463, 2031.25261020742, 1913.43246765846, 
    1796.92732439317, 1657.65058917257,
  4936.26514584792, 4123.6357475341, 3377.20733284678, 2889.1957547043, 
    2565.72896416456, 2288.40408515863, 2054.03968860635, 1922.30446863945, 
    1770.74787520852, 1663.55055916978,
  4959.91321608387, 4144.08787752412, 3329.15644996989, 2899.65840937701, 
    2513.33518797497, 2282.04684088801, 2058.73529740474, 1897.6959920311, 
    1761.52178717246, 1660.58321432322,
  4935.30173191977, 4197.71466212771, 3394.57516736225, 2867.3620031015, 
    2557.17972702811, 2250.3571611728, 2047.78290592795, 1896.29564319899, 
    1750.86184593294, 1665.22330403009 ;

 mean_source =
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000059, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000049, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000054, 0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000055, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.0000000000006, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000044, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000054, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000048, 0.10000000000005, 0.10000000000005, 0.10000000000005, 
    0.10000000000005, 0.10000000000005, 0.10000000000005, 0.10000000000005, 
    0.10000000000005, 0.10000000000005,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000038, 0.100000000000039, 0.100000000000039, 0.100000000000039, 
    0.100000000000039, 0.100000000000039, 0.100000000000039, 
    0.100000000000039, 0.100000000000039, 0.100000000000039,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000045, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000037, 0.100000000000038, 0.100000000000038, 0.100000000000038, 
    0.100000000000038, 0.100000000000038, 0.100000000000038, 
    0.100000000000038, 0.100000000000038, 0.100000000000038,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000047, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000054, 0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.0000000000003, 0.100000000000032, 0.100000000000032, 0.100000000000032, 
    0.100000000000032, 0.100000000000032, 0.100000000000032, 
    0.100000000000032, 0.100000000000032, 0.100000000000032,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.00000000000029, 0.10000000000003, 0.10000000000003, 0.10000000000003, 
    0.10000000000003, 0.10000000000003, 0.10000000000003, 0.10000000000003, 
    0.10000000000003, 0.10000000000003,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000056, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000052, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000043, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000063, 0.100000000000064, 0.100000000000064, 0.100000000000064, 
    0.100000000000064, 0.100000000000064, 0.100000000000064, 
    0.100000000000064, 0.100000000000064, 0.100000000000064,
  1.00000000000044, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000046, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000043, 0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000069, 0.10000000000007, 0.10000000000007, 0.10000000000007, 
    0.10000000000007, 0.10000000000007, 0.10000000000007, 0.10000000000007, 
    0.10000000000007, 0.10000000000007,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000055, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000062, 0.100000000000063, 0.100000000000063, 0.100000000000063, 
    0.100000000000063, 0.100000000000063, 0.100000000000063, 
    0.100000000000063, 0.100000000000063, 0.100000000000063,
  1.00000000000035, 0.100000000000036, 0.100000000000036, 0.100000000000036, 
    0.100000000000036, 0.100000000000036, 0.100000000000036, 
    0.100000000000036, 0.100000000000036, 0.100000000000036,
  1.00000000000049, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.00000000000035, 0.100000000000037, 0.100000000000037, 0.100000000000037, 
    0.100000000000037, 0.100000000000037, 0.100000000000037, 
    0.100000000000037, 0.100000000000037, 0.100000000000037,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000047, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000047, 0.100000000000048, 0.100000000000048, 0.100000000000048, 
    0.100000000000048, 0.100000000000048, 0.100000000000048, 
    0.100000000000048, 0.100000000000048, 0.100000000000048,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000058, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006,
  1.00000000000043, 0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044 ;

 source =
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000059, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000049, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000054, 0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000055, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.0000000000006, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000044, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000054, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000048, 0.10000000000005, 0.10000000000005, 0.10000000000005, 
    0.10000000000005, 0.10000000000005, 0.10000000000005, 0.10000000000005, 
    0.10000000000005, 0.10000000000005,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000038, 0.100000000000039, 0.100000000000039, 0.100000000000039, 
    0.100000000000039, 0.100000000000039, 0.100000000000039, 
    0.100000000000039, 0.100000000000039, 0.100000000000039,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000045, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000037, 0.100000000000038, 0.100000000000038, 0.100000000000038, 
    0.100000000000038, 0.100000000000038, 0.100000000000038, 
    0.100000000000038, 0.100000000000038, 0.100000000000038,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000047, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000054, 0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055, 
    0.100000000000055, 0.100000000000055, 0.100000000000055,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.0000000000003, 0.100000000000032, 0.100000000000032, 0.100000000000032, 
    0.100000000000032, 0.100000000000032, 0.100000000000032, 
    0.100000000000032, 0.100000000000032, 0.100000000000032,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.00000000000029, 0.10000000000003, 0.10000000000003, 0.10000000000003, 
    0.10000000000003, 0.10000000000003, 0.10000000000003, 0.10000000000003, 
    0.10000000000003, 0.10000000000003,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000046, 0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047, 
    0.100000000000047, 0.100000000000047, 0.100000000000047,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.0000000000006, 0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061, 
    0.100000000000061, 0.100000000000061, 0.100000000000061,
  1.00000000000056, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000052, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000043, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000063, 0.100000000000064, 0.100000000000064, 0.100000000000064, 
    0.100000000000064, 0.100000000000064, 0.100000000000064, 
    0.100000000000064, 0.100000000000064, 0.100000000000064,
  1.00000000000044, 0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045, 
    0.100000000000045, 0.100000000000045, 0.100000000000045,
  1.00000000000046, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000053, 0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054, 
    0.100000000000054, 0.100000000000054, 0.100000000000054,
  1.00000000000043, 0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000069, 0.10000000000007, 0.10000000000007, 0.10000000000007, 
    0.10000000000007, 0.10000000000007, 0.10000000000007, 0.10000000000007, 
    0.10000000000007, 0.10000000000007,
  1.00000000000057, 0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058, 
    0.100000000000058, 0.100000000000058, 0.100000000000058,
  1.00000000000055, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000048, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000051, 0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052, 
    0.100000000000052, 0.100000000000052, 0.100000000000052,
  1.00000000000062, 0.100000000000063, 0.100000000000063, 0.100000000000063, 
    0.100000000000063, 0.100000000000063, 0.100000000000063, 
    0.100000000000063, 0.100000000000063, 0.100000000000063,
  1.00000000000035, 0.100000000000036, 0.100000000000036, 0.100000000000036, 
    0.100000000000036, 0.100000000000036, 0.100000000000036, 
    0.100000000000036, 0.100000000000036, 0.100000000000036,
  1.00000000000049, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.00000000000055, 0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056, 
    0.100000000000056, 0.100000000000056, 0.100000000000056,
  1.00000000000056, 0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057, 
    0.100000000000057, 0.100000000000057, 0.100000000000057,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.00000000000035, 0.100000000000037, 0.100000000000037, 0.100000000000037, 
    0.100000000000037, 0.100000000000037, 0.100000000000037, 
    0.100000000000037, 0.100000000000037, 0.100000000000037,
  1.00000000000061, 0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062, 
    0.100000000000062, 0.100000000000062, 0.100000000000062,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.00000000000047, 0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049, 
    0.100000000000049, 0.100000000000049, 0.100000000000049,
  1.00000000000047, 0.100000000000048, 0.100000000000048, 0.100000000000048, 
    0.100000000000048, 0.100000000000048, 0.100000000000048, 
    0.100000000000048, 0.100000000000048, 0.100000000000048,
  1.00000000000045, 0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046, 
    0.100000000000046, 0.100000000000046, 0.100000000000046,
  1.0000000000004, 0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041, 
    0.100000000000041, 0.100000000000041, 0.100000000000041,
  1.0000000000005, 0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051, 
    0.100000000000051, 0.100000000000051, 0.100000000000051,
  1.00000000000052, 0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053, 
    0.100000000000053, 0.100000000000053, 0.100000000000053,
  1.00000000000058, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006, 0.10000000000006, 0.10000000000006, 
    0.10000000000006, 0.10000000000006,
  1.00000000000043, 0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044, 
    0.100000000000044, 0.100000000000044, 0.100000000000044 ;

 source_phase =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wind =
  19.6249309700917, 21.5090663232168, 21.7106667483167, 20.9468577089314, 
    23.0131307612275, 28.1839652464673, 22.6414755008295, 19.4443073967755, 
    22.3984046305349, 19.2968102953091,
  22.2316655347344, 20.5427104589286, 17.9117516231473, 18.7697229955621, 
    22.8316428674858, 25.7143543474726, 21.9545913336934, 24.8067374951338, 
    23.0788890663958, 22.3194100973918,
  20.5059989883605, 18.8306649090816, 20.1775464716551, 22.2439684567796, 
    19.083630303592, 18.9790795900592, 22.0374711383551, 22.9326508867602, 
    24.4288433821659, 21.9880803185923,
  17.1724512128409, 17.305157571735, 19.7920244207332, 20.0069290891, 
    24.3515590995139, 22.5804825546755, 18.3106449495295, 18.6753455130594, 
    20.1270350853068, 19.056631379356,
  23.019351041962, 23.480901556962, 20.8555915757753, 21.9748037892347, 
    26.9665259939397, 23.8471099345118, 25.2861039271466, 22.0343804070351, 
    22.3924082278445, 19.8392357484607,
  20.2367295992554, 19.4982257706854, 17.329340214301, 20.2345187885489, 
    23.8090784799045, 22.6517593379766, 18.8078528130198, 20.5890415127316, 
    23.3933454187276, 19.4087892823654,
  20.5167746059388, 19.8500562169152, 20.6982217550196, 23.6163283684632, 
    24.9312177652109, 24.462451798162, 21.8215964366857, 22.3179028060486, 
    24.2383307722412, 21.9623416907229,
  21.350150479496, 20.1893759882079, 19.753874828048, 18.7795239204614, 
    25.1839081852941, 25.6438817183165, 20.7572219386085, 21.8155187814719, 
    23.1732997058887, 22.3611640647658,
  19.4118601903101, 21.8460783620366, 21.1796923440267, 20.3351976280722, 
    22.2496413285256, 25.4278807509192, 22.4377425681452, 24.3206838548164, 
    22.0577708637598, 23.3010774047001,
  19.1611434651882, 18.4344524047594, 18.7152968720742, 18.1101381675083, 
    23.8487664243109, 23.8977178072767, 19.7823589299387, 21.2594144445519, 
    22.4490267547648, 21.6847467869033,
  21.2110029195181, 17.6484884388507, 19.2673152827467, 21.7801699316543, 
    24.1547831891127, 22.4032029916848, 21.464146386741, 21.5033623110365, 
    20.3441245841852, 22.2676649364405,
  18.2771565495209, 19.1977587890325, 17.370185283154, 20.3760920427319, 
    23.86616739763, 21.1014372731159, 17.6676703353542, 21.930008066689, 
    23.4657124540899, 20.9604557321403,
  18.555251626707, 20.3122700705233, 20.4013724494864, 18.6303968095356, 
    22.5603611768601, 23.7360813881301, 21.6472565551653, 21.716840919151, 
    22.7660361896531, 21.2234333565076,
  20.6703244747845, 16.800654079263, 19.0883021337656, 19.882702899903, 
    22.4000983052207, 23.2139122361521, 22.5651718641912, 21.4732079107684, 
    18.5697287632558, 19.5568925610897,
  19.8730455604997, 20.9920530569556, 21.5828093996238, 22.7257482677516, 
    25.4476652646715, 24.57793994888, 23.3779200122806, 21.250804544983, 
    22.4233924882603, 22.3163670884164,
  22.4546914515533, 21.8925564067937, 20.7883653395199, 25.2726980472426, 
    26.3039670335987, 23.142683711071, 19.9159138308777, 22.3041184623659, 
    23.1663507024909, 23.618691314097,
  17.3170429141094, 18.5621938381243, 17.6108980596626, 19.712813751723, 
    24.4074391188448, 21.8980223222239, 21.4141152146122, 19.7026610938911, 
    17.6648236332301, 20.2679647319594,
  20.4335450043158, 19.322099996281, 19.7061147342422, 19.7156067162985, 
    20.3229287133707, 26.7421134469238, 18.2389383483307, 21.8441941272217, 
    17.5820490755836, 24.4393629954678,
  22.008962824118, 20.3099201923761, 20.9255141828193, 22.2228389084524, 
    22.5715864693612, 22.4653404207663, 20.0582679043621, 20.6667265056376, 
    21.5616710711408, 22.42263233972,
  19.3354636279061, 20.7230826642697, 19.2475274788118, 20.8278417989833, 
    22.8975338239968, 20.9819160760162, 21.0716164637633, 21.9767302256232, 
    18.7879530301013, 19.395587565909,
  18.7842223605985, 20.8361436500519, 22.2506947749683, 17.8263792860035, 
    20.3375429054526, 24.5990226112524, 20.7560045975247, 21.3276375560733, 
    22.9992765059053, 23.3032271577844,
  19.2163403746698, 20.107177866568, 20.6521801895324, 20.7391998564355, 
    24.0220721993147, 24.9082033590743, 23.0706465199116, 22.7134392699063, 
    21.0572912964982, 22.466146057007,
  21.585853690655, 20.566922232807, 20.9588170080915, 22.0647589441024, 
    25.5009587085965, 26.1014448370435, 21.6414764487554, 24.9246565912923, 
    25.3223558591914, 23.8516887940137,
  23.2701356940825, 22.2234611971093, 24.2012341138996, 23.7800804881245, 
    26.0074332943245, 26.5714291990976, 22.3668043093078, 26.8037111898027, 
    22.3063223073737, 23.9429436796466,
  21.3869505079468, 21.7129995660199, 21.1171899839701, 20.194956237949, 
    24.9072904220401, 23.218608675045, 24.1753051485497, 24.3708901259122, 
    23.8303716186174, 23.0685792808097,
  21.2139652903025, 18.4538943175751, 18.6621911950968, 20.7467528847222, 
    18.6581006837334, 25.2229918457611, 22.0511618407268, 20.8345137511958, 
    22.0497425340889, 18.3684068397101,
  20.1818621909498, 18.9098301253293, 22.0436960423488, 18.7670339281514, 
    26.2117801528981, 22.8385666736169, 21.6346989128121, 21.8853073302088, 
    19.9986955248676, 23.2749737741453,
  19.4661538913934, 17.5861619117166, 18.8635932072729, 19.7035433491066, 
    22.5783916519968, 23.6920786515433, 18.6267046665279, 22.4714271543035, 
    21.7722527105653, 18.9400925168309,
  20.1080538147119, 20.668094742738, 19.1541157724254, 18.7485333171167, 
    22.1620419503362, 23.5721533022712, 20.6005047304139, 19.5728200109686, 
    18.8442617927029, 21.8179675754862,
  20.9223522622115, 19.1121232672422, 20.1274643469491, 21.4287687868367, 
    26.5387087449504, 23.454942241408, 22.714543976311, 24.0447663919274, 
    23.4413436074889, 20.1498678378216,
  19.3769990574516, 19.3470251641666, 19.2021207283676, 18.019037822923, 
    25.1744498065142, 22.6823781780647, 21.9127776381343, 17.4540100866893, 
    20.6708559988149, 22.3543376949761,
  19.3670644064467, 19.1076703604091, 18.8854808802279, 20.7416009664874, 
    20.2718675760211, 24.875141955296, 19.2554601628667, 19.3126868688605, 
    22.3122158955327, 20.731784848084,
  19.7749589309895, 20.9144362131247, 22.4435782192791, 22.7471279374615, 
    23.8131758092616, 26.2274332381142, 22.4553568383611, 21.2496467968501, 
    22.423368177464, 23.5686062310841,
  20.3939618381091, 20.0787711286317, 20.7771909178821, 22.6507888659002, 
    22.8313974551788, 26.2517383517316, 22.5669763608782, 22.5565518774206, 
    22.4917816304608, 22.6018870913256,
  23.5189606818689, 19.0294794788023, 20.7160207935934, 22.2834460844027, 
    21.4194477049157, 26.3137917903553, 23.642464010342, 22.9152253504596, 
    20.697755896371, 25.0739256832045,
  17.7726189475035, 20.0081163320631, 20.0458298079193, 22.3066833694154, 
    22.8221026861796, 27.5558561638423, 22.7656481257465, 23.9815370934922, 
    22.7415097553971, 20.0498836817772,
  19.4269394591382, 19.8061223956145, 18.7633293912859, 19.3703330512199, 
    23.3378142832975, 23.6304028857352, 23.1161444296917, 20.0717248659881, 
    19.732052540028, 21.0734765001828,
  20.8770746127703, 19.5267849827676, 19.0781590495218, 21.2731172061216, 
    22.4237253904994, 22.5733209975188, 20.877855362113, 22.7386521192746, 
    24.5367133212109, 21.3198289313593,
  19.4960998279283, 19.7271240973046, 16.8906283524408, 17.5750207785723, 
    22.6974529686628, 23.6310912756864, 20.7588536330908, 20.5618925266947, 
    19.4939581585775, 22.0083059859112,
  18.1867495314236, 19.3170618155341, 19.7846396523151, 22.9349558868561, 
    25.729708621553, 27.4951850795233, 23.2208095773663, 23.3654065411441, 
    21.8337768531952, 18.3243807865392,
  22.2582569771423, 21.6073946758329, 21.7043560959378, 23.3745948625747, 
    26.4942274533129, 26.733752077764, 23.8648983986641, 23.2608542850248, 
    24.1121053081357, 20.180701686042,
  21.4566428265671, 18.5394135283347, 17.6657357527022, 19.0628236639948, 
    22.7447084956596, 22.0160200822911, 20.957773540365, 22.6761319127668, 
    18.9836864369893, 18.5087088899513,
  22.944503543479, 21.0155090762187, 18.5338342524752, 23.0329918781166, 
    24.4223893567573, 24.0665586281184, 21.3155514475258, 24.4875568290283, 
    25.178902207332, 21.026928164455,
  21.8139918738416, 20.6721848656404, 19.5296416108205, 21.8688563512069, 
    24.3327266555838, 23.1723790327946, 20.587018709315, 19.0984696300328, 
    21.3461475944063, 24.0878366197193,
  21.9978595628748, 20.1504385092186, 21.4166615130902, 21.2576936113091, 
    25.6910499036806, 23.1794011966747, 24.3584276454134, 23.8024455696118, 
    24.2492370872677, 24.6914583414172,
  16.5904444085935, 17.6257325771034, 18.2551546681909, 20.2099426336598, 
    21.609140059341, 21.5335288507248, 19.5613578277287, 20.5120964767494, 
    19.7931216423593, 19.3789846809258,
  20.1845417047926, 18.3727504162256, 20.8640132798357, 18.8688759343258, 
    22.0137199531165, 24.2050326767379, 19.8108593606415, 17.8063992006127, 
    23.2633409343208, 21.4861463087443,
  19.6518729286276, 20.2388925745753, 22.5530430682637, 22.7784719025498, 
    24.8570957659204, 26.2528576191955, 22.3864112165413, 24.2599488147884, 
    22.2678561920121, 21.5942313115748,
  20.1907764004336, 19.5147981731442, 21.2624568157203, 20.3950068112795, 
    22.656077657414, 24.2680639548654, 22.5526260529477, 21.8338703731042, 
    22.5313077920591, 22.2631691379656,
  21.1643653568738, 19.8826965558811, 20.2275705213433, 20.0021132626311, 
    23.3158753912755, 23.6047282178929, 25.6287949479375, 23.1510390117148, 
    23.21924229509, 21.882033400218,
  22.1460663281232, 20.2390152489265, 19.039374327701, 19.7666314355337, 
    26.1403065056624, 26.7959784400582, 21.3414506625264, 21.446176289424, 
    22.4345946044741, 22.2986460948746,
  19.240375279715, 20.6659838374038, 19.2866566643194, 20.1002730614372, 
    26.000519261987, 24.0408313490448, 22.6531235388352, 22.0477040122371, 
    22.882746612423, 20.0926905691669,
  20.3520908633866, 19.9086714792572, 20.3559190450373, 19.6060500528339, 
    26.2630425870344, 24.6833533587566, 20.3319347552104, 20.2074694929196, 
    21.2001353248893, 22.4151748276326,
  21.176837448357, 17.5867033334996, 17.7030050694566, 20.7350537802925, 
    22.4288354412503, 23.0306891666961, 19.1178436111304, 20.699555393153, 
    19.7960300147495, 18.6564598616604,
  20.044274898024, 20.3669632715759, 17.9343174092219, 19.7687801828674, 
    22.9049357388899, 23.3278475041481, 21.4632669178636, 22.2908112619707, 
    21.0803173434389, 21.4932088957938,
  21.6062375929694, 22.5236622667373, 20.0733896226814, 19.8918055526762, 
    23.0969102876787, 23.2058855192561, 19.4780787697965, 21.984180810592, 
    21.1912025077916, 21.8426285765593,
  22.1343430708991, 19.9136070594121, 20.7320407397566, 21.364775149414, 
    23.4013410680772, 22.1116479312564, 20.0344828852105, 21.9018916991106, 
    21.6614156241361, 20.5616102217979,
  21.9827603208728, 20.7530414297835, 16.7802646613637, 22.2895627401528, 
    23.6399601138275, 23.6117352370409, 21.0795235173053, 23.2678265630638, 
    23.5156223706717, 23.1875665316692,
  20.493498409572, 21.8151151050499, 21.9066413427573, 22.8156949840686, 
    24.3679090954473, 23.4547500022643, 20.4451875921773, 20.6665825496724, 
    20.7502078948482, 21.8735038592288,
  20.3359820148419, 20.4629700028859, 18.0970616781538, 20.1572491614619, 
    23.0130975624218, 22.4328801563887, 20.8197288141429, 21.1839328344749, 
    22.2238283763054, 21.207249351023,
  20.6462610953227, 20.6043047405246, 19.6379242844012, 22.2019946621877, 
    23.4289777820152, 24.8265982529431, 20.4329398742808, 23.1859892208646, 
    24.2635303839843, 25.081854624701,
  22.0776842440405, 19.2013928120267, 19.8071569872927, 22.2201224340338, 
    26.5687051437968, 27.7192170161072, 22.705502202708, 23.4747365660503, 
    21.4665986090492, 23.0594067034969,
  20.2925691863507, 17.7751668909402, 18.4039047238961, 16.7631838617413, 
    21.2879114124662, 23.6696001936749, 19.6075592992575, 20.624669149067, 
    21.6524285323945, 19.7819934282455,
  18.1054158426523, 19.9989102219346, 20.7834909563412, 18.9665278707828, 
    25.4854205973084, 24.4426613505103, 22.5325971005892, 24.1827277090218, 
    21.4832859688028, 23.5964743490822,
  22.6752343097278, 19.9502636611785, 18.2391452471715, 21.1030814924503, 
    21.9559150655741, 24.1558314972333, 19.9305249401331, 25.4022140317211, 
    21.2933606035308, 22.8797263379449,
  18.3548144272872, 19.9130910486747, 18.7439002539931, 23.4647939986876, 
    23.9435983660278, 26.1881134544215, 21.3295389760177, 22.2057989321621, 
    24.2265432000508, 23.0300808264806,
  21.9856550930253, 18.8099678156943, 17.4752128803057, 20.3136839352391, 
    21.1430442537274, 21.8911468648469, 22.2235402755766, 23.5544499121218, 
    19.9327967802021, 22.0884227902946,
  20.8039737800154, 18.5491165739058, 19.8483570238978, 19.6577586334409, 
    22.7293019186313, 27.3669535429267, 23.6722506398789, 21.9876495909018, 
    23.5934751960555, 22.4336911574151,
  19.0215049348978, 18.6244911813375, 18.1543003542628, 20.8386454028469, 
    23.6350563426476, 22.5284662433271, 22.8332651514022, 22.8260856383512, 
    24.3001306386811, 22.6273281670919,
  22.284914067416, 20.4786678851048, 18.5699150486217, 19.9723896798977, 
    24.8894646863479, 24.0577296926846, 18.716992004327, 24.4897548093821, 
    22.3318635141275, 23.7708474318921,
  21.8260070656087, 22.4097846730676, 18.4702606029232, 21.2037674357942, 
    26.49667674596, 25.893941723468, 23.3603225903716, 23.9075204008819, 
    20.3596525390173, 24.2972555162252,
  21.5573715729374, 21.1612522626769, 22.3758802358839, 21.4469974655204, 
    25.2981380680944, 24.2145960808384, 21.757962082981, 23.1597171259488, 
    24.5787533282042, 23.1470641744999,
  18.3974057083314, 18.6780544941245, 18.0807000809553, 18.5325666428358, 
    23.3327722261678, 21.4738912243292, 20.9990125362725, 20.0078199993289, 
    18.3832367524686, 18.8023609848967,
  21.9491810525246, 19.7716779544379, 18.5465509500256, 20.3072882816021, 
    23.5731400948066, 22.9144415582392, 19.0759823467407, 23.8478638181577, 
    23.7168975482792, 20.4389762614991,
  18.9361913560642, 21.0946871871436, 21.2300887557843, 21.5800524811259, 
    21.3056008863743, 24.8274853057091, 21.1328400356026, 21.5548638612101, 
    23.7355312871334, 21.1991623942634,
  21.4774632555289, 18.9169585399884, 20.6874722548899, 21.5853500736947, 
    23.112433973902, 23.445946959647, 20.2327258710806, 20.8240453009503, 
    21.4981566663487, 21.4608473203805,
  18.0315710878689, 21.5372152964458, 19.4193572259521, 20.3444777976534, 
    25.2730366548758, 26.2927741043476, 20.4759068646439, 22.3123500931917, 
    24.4671848848749, 22.7776968357497,
  20.6636975967031, 20.355040953058, 19.6383845756746, 20.5558926165957, 
    25.2420359879901, 23.6702712853034, 23.8391577224089, 22.0939907173268, 
    21.9456945517534, 22.0665616114532,
  21.3248985367175, 19.2315682429829, 18.4616805190862, 19.0238352645292, 
    23.8376714285204, 22.2766779513412, 22.2101662076882, 24.5233219471702, 
    21.860996187177, 20.3668661693499,
  21.4058803998674, 19.2040592980853, 21.311536146935, 23.7417488540893, 
    24.287964568376, 23.801229879017, 18.3383516539401, 22.5385628386695, 
    21.3148663946344, 19.6583711575979 ;

 concentration_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mean_source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_phase_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wind_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 concentration_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 mean_source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_phase_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 wind_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 location = 0, 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9 ;

 time = 41.666666666666667 ;

 advance_to_time = 41.666666666666667 ;
}
