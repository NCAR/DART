netcdf wrf_input {
dimensions:
	Times = 37 ;
	x = 3 ;
	y = 3 ;
	x_stag = 4 ;
	y_stag = 4 ;
	z_amsl = 34 ;
	z_amsl_stag = 35 ;
	variable_scr = 4 ;
	variable_sfc = 11 ;
	soil_levels = 4 ;
	variable_soil = 2 ;
	ext_scalar = 1 ;
	record = UNLIMITED ; 
variables:
	int inityear(record, Times) ;
	int initmonth(record, Times) ;
	int initday(record, Times) ;
	int inithour(record, Times) ;
	float Z(record, Times, z_amsl_stag, y, x) ;
	float T(record, Times, z_amsl, y, x) ;
		T:_FillValue = -999.f ;
	float Q(record, Times, z_amsl, y, x) ;
	float P(record, Times, z_amsl, y, x) ;
	float U(record, Times, z_amsl, y, x_stag) ;
	float V(record, Times, z_amsl, y_stag, x) ;
	float PRECIP(record, Times, y, x) ;
	float MU(record, Times, y, x) ;
	float MUB(record, Times, y, x) ;
	float MU0(record, Times, y, x) ;
	float ZNU(record, Times, z_amsl) ;
	float ZNW(record, Times, z_amsl_stag) ;
	float P_TOP(record, Times, ext_scalar) ;
	float MAPFAC_M(record, Times, y, x) ;
	float screen(record, Times, y, x, variable_scr) ;
		screen:_FillValue = -999.f ;
	float surface(record, Times, y, x, variable_sfc) ;
		surface:_FillValue = -999.f ;
	float soil(record, Times, soil_levels, y, x, variable_soil) ;
		soil:_FillValue = -999.f ;
	float lats(record, Times, y, x) ;
	float lons(record, Times, y, x) ;
	float terrain(record, Times, y, x) ;

// global attributes:
		:misc_order = "PBLH" ;
		:soil_order = "TSLB,SMOIS" ;
		:sfc_order = "TSK,GLW,GSW,TMN,HFX,QFX,QSFC,VEGFRA,ISLTYP,IVGTYP,LU_INDEX" ;
		:screen_order = "T2,U10,V10,Q2(mixing ratio)" ;
		:times = "4-hourly" ;
		:contents = "profiles from WRF 4KM BAMEX run" ;
		:creation_date = "Mon Dec 19 22:06:27 MST 2005" ;
		:TITLE = " OUTPUT FROM WRF V1.3 MODEL" ;
		:START_DATE = "2003-05-03_00:00:00" ;
		:WEST-EAST_GRID_DIMENSION = 501 ;
		:SOUTH-NORTH_GRID_DIMENSION = 501 ;
		:BOTTOM-TOP_GRID_DIMENSION = 34 ;
		:DYN_OPT = 2 ;
		:DIFF_OPT = 1 ;
		:KM_OPT = 4 ;
		:DAMP_OPT = 0 ;
		:KHDIF = 0.f ;
		:KVDIF = 0.f ;
		:MP_PHYSICS = 2 ;
		:RA_LW_PHYSICS = 1 ;
		:RA_SW_PHYSICS = 1 ;
		:BL_SFCLAY_PHYSICS = 1 ;
		:BL_SURFACE_PHYSICS = 2 ;
		:BL_PBL_PHYSICS = 1 ;
		:CU_PHYSICS = 0 ;
		:WEST-EAST_PATCH_START_UNSTAG = 377 ;
		:WEST-EAST_PATCH_END_UNSTAG = 500 ;
		:WEST-EAST_PATCH_START_STAG = 377 ;
		:WEST-EAST_PATCH_END_STAG = 501 ;
		:SOUTH-NORTH_PATCH_START_UNSTAG = 485 ;
		:SOUTH-NORTH_PATCH_END_UNSTAG = 500 ;
		:SOUTH-NORTH_PATCH_START_STAG = 485 ;
		:SOUTH-NORTH_PATCH_END_STAG = 501 ;
		:BOTTOM-TOP_PATCH_START_UNSTAG = 1 ;
		:BOTTOM-TOP_PATCH_END_UNSTAG = 34 ;
		:BOTTOM-TOP_PATCH_START_STAG = 1 ;
		:BOTTOM-TOP_PATCH_END_STAG = 35 ;
		:DX = 4000.f ;
		:DY = 4000.f ;
		:DT = 24.f ;
		:CEN_LAT = 40.00001f ;
		:CEN_LON = -95.f ;
		:TRUELAT1 = 30.f ;
		:TRUELAT2 = 45.f ;
		:GMT = 0.f ;
		:JULYR = 2003 ;
		:JULDAY = 123 ;
		:ISWATER = 16 ;
		:MAP_PROJ = 1 ;
		:MMINLU = "USGS" ;
		:SW_LON = -105.4442f ;
		:SW_LAT = 30.46228f ;
}
