netcdf sondes_obs_2018041500.200 {
dimensions:
	Location = 200 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 974LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:date_time = 2018041500 ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
		:history = "Tue Jul 22 15:18:20 2025: ncks -dLocation,0,199 IODA_READERS/UKMO/INPUTS/sondes_obs_2018041500_m.nc4 sondes_obs_2018041500_m.200.nc4\nWed Apr 10 16:32:50 2024: ncrename -v .sensorChannelNumber,Channel ./sondes_obs_2018041500_m.nc4 ./data2/sondes_obs_2018041500_m.nc4\nWed Nov 23 02:47:22 2022: ncks --cnk_dmn Location,100 -L 4 new.nc4 sondes_obs_2018041500_m.nc4" ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

group: GsiAdjustObsError {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  data:

   airTemperature = _, _, 1.024938, _, _, 1.139351, _, 1.534971, 1.051251, _, 
      1.050533, 1.401237, _, _, 1.2, _, 1.145388, _, _, _, 1.68, _, _, _, 
      0.96, _, _, _, _, _, 1.29849, 2.122585, _, 2.12298, 1.294087, _, _, 
      1.314831, _, 1.32547, _, _, 1.08, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, 1.8, 1.8, _, 1.8, 1.68, 1.68, 1.32, 1.08, 1.8, 
      1.8, 0.96, 1.56, 1.2, 1.08, 1, 1.212887, 1.2, 0.96, 1.41979, 1.931882, 
      1.448028, 0.8, 1, _, 1.1, 1.343928, 1.343936, 1.2, 1.2, 1.1, 1, 
      0.9872137, 0.9848667, 0.96, 1.08, 1.2, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, 0.96, 1.2, 1.08, 0.8, 1.2, 1.44, 2.12298, 
      2.122585, 1.56, 1.56, 1.8, 1.8, 1.8, 1, 1.626305, 1.626304, 1.2, 1, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 10.56813, 9.957422, 10.09526, 11.06756, 
      12.00879, 16.53376, 23.17653, 35.09987, 8.544992e-05, 0.0001147122, 
      0.0001975877, 0.0002286237, 0.0003814484, _, 0.0009811161, 
      0.0009813248, 0.0004945507, 0.0009753293, 0.0008994794, 0.0005680757, 
      0.0006505361, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      14.31543, 11.10419, 10.03266, 24.07659, 9.466661, 23.28926, 19.19881, 
      22.04181, 5.867995, 21.62867, 31.04534, 8.654429, 5.022742, 6.947986, 
      12.853, 54.1556, 7.45339, 11.96863, 0.003287753, 43.96388, 8.303241, 
      7.985352, 0.003925482, 63.1524, 0.004738071, 5.541402, 0.006204558, 
      0.008775169, 0.005110189, 6.162792, 5.046216, 111.7017, 106.5203, 
      66.78051, 4.642167, 184.0855, 87.48625, 0.0002088464, 99.78229, 
      0.0002302065, 0.0002566602, 0.00042202, 0.0005839344, 0.001844437, 
      0.0009510599, 0.0008013952, 0.0005883959, 0.0008268948, 0.0007247257, 
      0.001465403, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 2.3, 2.933219, _, 2.933222, 2.269284, _, 2.513141, _, _, 
      2.441647, _, _, 2.5, 3.795623, _, 3.248051, _, 3.598207, 3.191818, 2.1, 
      _, 2.52, 2.1, 2.1, _, 2.52, 2.1, 2.105534, 2.52, 2.254568, _, _, 2.52, 
      _, _, 2.678262, 2.52, _, 2.52, _, 3.1, 2.52, _, 3.229246, 1.59254, _, 
      1.590933, 1.4, 1.5, 1.5, 3.975462, 3.989056, 1.659325, 1.651189, 1.6, 
      3.101022, 3.101012, 1.6, 1.6, 2.337516, 2.337529, 1.9, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      2.195697, 2.7, 2.9, 3.1, 3.66084, 5.976196, 4.755991, 3.214425, 
      3.627078, 3.627078, 2.9, 2.8, 2.924455 ;

   windNorthward = 2.3, 2.933219, _, 2.933222, 2.269284, _, 2.513141, _, _, 
      2.441647, _, _, 2.5, 3.795623, _, 3.248051, _, 3.598207, 3.191818, 2.1, 
      _, 2.52, 2.1, 2.1, _, 2.52, 2.1, 2.105534, 2.52, 2.254568, _, _, 2.52, 
      _, _, 2.678262, 2.52, _, 2.52, _, 3.1, 2.52, _, 3.229246, 1.59254, _, 
      1.590933, 1.4, 1.5, 1.5, 3.975462, 3.989056, 1.659325, 1.651189, 1.6, 
      3.101022, 3.101012, 1.6, 1.6, 2.337516, 2.337529, 1.9, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      2.195697, 2.7, 2.9, 3.1, 3.66084, 5.976196, 4.755991, 3.214425, 
      3.627078, 3.627078, 2.9, 2.8, 2.924455 ;
  } // group GsiAdjustObsError

group: GsiFinalObsError {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  data:

   airTemperature = _, _, 1.024938, _, _, 1.139351, _, 1.534971, 1.051251, _, 
      1.050533, 1.401237, _, _, 1.2, _, 1.145388, _, _, _, 1.68, _, _, _, 
      0.96, _, _, _, _, _, 1.29849, 2.122585, _, 2.12298, 1.294087, _, _, 
      1.314831, _, 1.32547, _, _, 1.08, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, 1.8, 1.8, _, 1.8, 1.68, 1.68, 1.32, 1.08, 1.8, 
      1.8, 0.96, 1.56, 1.2, 1.08, 1, 1.212887, 1.2, 0.96, 1.41979, 1.931882, 
      1.448028, 0.8, 1, _, 1.1, 1.343928, 1.343936, 1.2, 1.2, 1.1, 1, 
      0.9872137, 0.9848667, 0.96, 1.08, 1.2, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, 0.96, 1.2, 1.08, 0.8, 1.2, 1.44, 2.12298, 
      2.122585, 1.56, 1.56, 1.8, 1.8, 1.8, 1, 1.626305, 1.626304, 1.2, 1, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 10.56813, 9.957422, 10.09526, 11.06756, 
      12.00879, 16.53376, 23.17653, 35.09987, 0.0001, 0.0001147122, 
      0.0001975877, 0.0002286237, 0.0003814484, _, 17.29257, 0.7433912, 
      0.0004945507, 0.0009753293, 0.0008994794, 0.0005680757, 0.0006505361, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 14.31543, 
      11.10419, 10.03266, 24.07659, 9.466661, 23.28926, 19.19881, 22.04181, 
      5.867995, 21.62867, 31.04534, 8.654429, 5.022742, 6.947986, 12.853, 
      54.1556, 7.45339, 11.96863, 0.003287753, 43.96388, 8.303241, 7.985352, 
      0.003925482, 63.1524, 0.004738071, 5.541402, 0.006204558, 6.511775, 
      9.486762, 6.162792, 5.046216, 111.7017, 106.5203, 66.78051, 4.642167, 
      184.0855, 87.48625, 0.0002088464, 99.78229, 0.0002302065, 0.0002566602, 
      0.00042202, 0.0005839344, 0.001844437, 0.0009510599, 0.0008013952, 
      0.0005883959, 0.0008268948, 0.0007247257, 0.001465403, _, _, _, _, _, 
      _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 100.0536, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      258.6004, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      178.2108, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 187.0397, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 2.3, 2.933219, _, 2.933222, 2.269284, _, 2.513141, _, _, 
      2.441647, _, _, 2.5, 3.795623, _, 3.248051, _, 3.598207, 3.191818, 2.1, 
      _, 2.52, 2.1, 2.1, _, 2.52, 2.1, 2.105534, 2.52, 2.254568, _, _, 2.52, 
      _, _, 2.678262, 2.52, _, 2.52, _, 3.1, 2.52, _, 3.229246, 1.671352, _, 
      1.590933, 1.4, 1.5, 1.5, 3.975462, 3.989056, 1.659325, 1.651189, 1.6, 
      3.101022, 3.101012, 1.6, 1.6, 2.337516, 2.337529, 1.9, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      2.195697, 2.7, 2.9, 3.1, 3.66084, 5.976196, 4.755991, 3.214425, 
      3.627078, 3.627078, 2.9, 2.8, 2.924455 ;

   windNorthward = 2.3, 2.933219, _, 2.933222, 2.269284, _, 2.513141, _, _, 
      2.441647, _, _, 2.5, 3.795623, _, 3.248051, _, 3.598207, 3.191818, 2.1, 
      _, 2.52, 2.1, 2.1, _, 2.52, 2.1, 2.105534, 2.52, 2.254568, _, _, 2.52, 
      _, _, 2.678262, 2.52, _, 2.52, _, 3.1, 2.52, _, 3.229246, 1.671352, _, 
      1.590933, 1.4, 1.5, 1.5, 3.975462, 3.989056, 1.659325, 1.651189, 1.6, 
      3.101022, 3.101012, 1.6, 1.6, 2.337516, 2.337529, 1.9, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      2.195697, 2.7, 2.9, 3.1, 3.66084, 5.976196, 4.755991, 3.214425, 
      3.627078, 3.627078, 2.9, 2.8, 2.924455 ;
  } // group GsiFinalObsError

group: GsiHofX {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  		string airTemperature:units = "K" ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  		string specificHumidity:units = "1" ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  		string stationPressure:units = "Pa" ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  		string windEastward:units = "m s-1" ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  		string windNorthward:units = "m s-1" ;
  data:

   airTemperature = _, _, 217.8734, _, _, 217.0876, _, 215.5437, 215.816, _, 
      215.8251, 214.9051, _, _, 213.0954, _, 213.341, _, _, _, 218.4771, _, 
      _, _, 215.8257, _, _, _, _, _, 215.4191, 216.1662, _, 216.1376, 
      215.3677, _, _, 214.6395, _, 214.5411, _, _, 214.9398, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, 220.4012, 220.7459, _, 
      218.8324, 217.6263, 216.191, 211.6831, 212.6178, 228.9244, 227.2065, 
      213.5374, 212.888, 211.4368, 212.6485, 221.0848, 220.497, 220.5779, 
      213.2851, 220.5432, 220.5466, 220.5248, 216.095, 218.9233, _, 218.1157, 
      218.6098, 218.917, 220.1382, 222.3568, 222.8333, 222.9289, 221.1145, 
      221.0343, 220.6421, 219.5625, 218.73, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, 219.153, 217.5795, 218.5904, 220.1139, 
      218.5044, 220.7928, 221.7886, 221.8312, 222.267, 222.7007, 228.9026, 
      230.0084, 227.0155, 221.6562, 221.7667, 221.7365, 219.4576, 219.5215, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 1.261783e-05, 1.61458e-05, 1.923614e-05, 
      2.131738e-05, 2.333161e-05, 3.195423e-05, 4.488333e-05, 6.8583e-05, 
      0.0001737459, 0.0002314164, 0.0003142061, 0.0003059815, 0.0002820091, 
      _, 0.002293864, 0.00229393, 0.0004977643, 0.001810573, 0.001568854, 
      0.0007475786, 0.001156733, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, 3.955063e-06, 5.602848e-06, 6.865373e-06, 5.211112e-06, 
      7.935005e-06, 5.06659e-06, 4.535333e-06, 4.849369e-06, 3.590828e-06, 
      4.803433e-06, 5.577111e-06, 8.150771e-06, 2.94438e-06, 3.816171e-06, 
      4.526688e-06, 5.345446e-06, 5.09409e-06, 4.408481e-06, 0.004212357, 
      6.773343e-06, 7.229421e-06, 6.425549e-06, 0.004611935, 5.675943e-06, 
      0.004862144, 2.362684e-06, 0.00503738, 0.005036596, 0.005036283, 
      2.685049e-06, 2.341293e-06, 2.130789e-05, 1.827357e-05, 7.142411e-06, 
      2.560825e-06, 5.536221e-05, 9.537472e-06, 6.951868e-05, 1.436888e-05, 
      9.297661e-05, 0.0001597527, 0.001088456, 0.0014386, 0.00348485, 
      0.001627005, 0.001658239, 0.001924701, 0.002191405, 0.002213344, 
      0.003280398, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 101088.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      101447, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      98670.73, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 92450.84, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 6.152787, 10.2754, _, 11.21958, 5.261633, _, 4.536641, _, 
      _, 4.108237, _, _, 14.65928, 13.87475, _, 14.09263, _, 13.40247, 
      15.28347, 2.949898, _, 7.738989, 2.874058, 2.913944, _, 6.160647, 
      2.68786, 2.007444, 5.093765, 2.018525, _, _, 4.455017, _, _, 2.12737, 
      3.534173, _, 4.242957, _, 28.79542, 3.990478, _, 28.61979, -1.904203, 
      _, -3.527674, -3.145489, -1.640043, 0.1895263, 17.29115, 16.96097, 
      3.877544, 4.56585, 5.699979, 13.75763, 13.93032, 5.559056, 5.670705, 
      10.86785, 10.40997, 7.717412, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -1.225706, 11.69911, 
      13.06857, 14.05671, 14.53291, 14.48116, 14.47679, 14.39564, 14.87393, 
      14.7753, 13.68717, 11.97302, 9.113683 ;

   windNorthward = 2.380202, -1.089164, _, -1.794114, 2.936322, _, 2.991843, 
      _, _, 3.023115, _, _, -1.289333, -5.006013, _, -4.117733, _, -7.001625, 
      -8.685597, 3.64881, _, -2.802598, 4.037339, 3.779823, _, -2.583868, 
      3.388475, 2.828758, -2.67919, 2.65556, _, _, -2.773853, _, _, 2.491153, 
      -2.889902, _, -2.150659, _, -14.0447, 0.8029721, _, -12.92819, 
      1.643805, _, 4.388265, 6.986234, 6.684765, 6.673048, -7.191293, 
      -6.860639, 5.680958, 5.309257, 4.528631, -0.4637186, -0.1207601, 
      3.963976, 3.485844, -2.31085, -2.212005, 0.5185826, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      -0.8737034, 1.998885, 1.880142, 1.405234, 0.3026514, -0.5946224, 
      -0.6703909, -2.077407, -5.476562, -6.520739, -11.21046, -12.62324, 
      -9.750257 ;
  } // group GsiHofX

group: GsiHofXBc {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  		string airTemperature:units = "K" ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  		string specificHumidity:units = "1" ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  		string stationPressure:units = "Pa" ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  		string windEastward:units = "m s-1" ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  		string windNorthward:units = "m s-1" ;
  data:

   airTemperature = _, _, 217.8734, _, _, 217.0876, _, 215.5437, 215.816, _, 
      215.8251, 214.9051, _, _, 213.0954, _, 213.341, _, _, _, 218.4771, _, 
      _, _, 215.8257, _, _, _, _, _, 215.4191, 216.1662, _, 216.1376, 
      215.3677, _, _, 214.6395, _, 214.5411, _, _, 214.9398, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, 220.4012, 220.7459, _, 
      218.8324, 217.6263, 216.191, 211.6831, 212.6178, 228.9244, 227.2065, 
      213.5374, 212.888, 211.4368, 212.6485, 221.0848, 220.497, 220.5779, 
      213.2851, 220.5432, 220.5466, 220.5248, 216.095, 218.9233, _, 218.1157, 
      218.6098, 218.917, 220.1382, 222.3568, 222.8333, 222.9289, 221.1145, 
      221.0343, 220.6421, 219.5625, 218.73, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, 219.153, 217.5795, 218.5904, 220.1139, 
      218.5044, 220.7928, 221.7886, 221.8312, 222.267, 222.7007, 228.9026, 
      230.0084, 227.0155, 221.6562, 221.7667, 221.7365, 219.4576, 219.5215, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 1.261783e-05, 1.61458e-05, 1.923614e-05, 
      2.131738e-05, 2.333161e-05, 3.195423e-05, 4.488333e-05, 6.8583e-05, 
      0.0001737459, 0.0002314164, 0.0003142061, 0.0003059815, 0.0002820091, 
      _, 0.002293864, 0.00229393, 0.0004977643, 0.001810573, 0.001568854, 
      0.0007475786, 0.001156733, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, 3.955063e-06, 5.602848e-06, 6.865373e-06, 5.211112e-06, 
      7.935005e-06, 5.06659e-06, 4.535333e-06, 4.849369e-06, 3.590828e-06, 
      4.803433e-06, 5.577111e-06, 8.150771e-06, 2.94438e-06, 3.816171e-06, 
      4.526688e-06, 5.345446e-06, 5.09409e-06, 4.408481e-06, 0.004212357, 
      6.773343e-06, 7.229421e-06, 6.425549e-06, 0.004611935, 5.675943e-06, 
      0.004862144, 2.362684e-06, 0.00503738, 0.005036596, 0.005036283, 
      2.685049e-06, 2.341293e-06, 2.130789e-05, 1.827357e-05, 7.142411e-06, 
      2.560825e-06, 5.536221e-05, 9.537472e-06, 6.951868e-05, 1.436888e-05, 
      9.297661e-05, 0.0001597527, 0.001088456, 0.0014386, 0.00348485, 
      0.001627005, 0.001658239, 0.001924701, 0.002191405, 0.002213344, 
      0.003280398, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 101045.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      101936.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      99714.68, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 93558.94, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 6.152787, 10.2754, _, 11.21958, 5.261633, _, 4.536641, _, 
      _, 4.108237, _, _, 14.65928, 13.87475, _, 14.09263, _, 13.40247, 
      15.28347, 2.949898, _, 7.738989, 2.874058, 2.913944, _, 6.160647, 
      2.68786, 2.007444, 5.093765, 2.018525, _, _, 4.455017, _, _, 2.12737, 
      3.534173, _, 4.242957, _, 28.79542, 3.990478, _, 28.61979, -1.904203, 
      _, -3.527674, -3.145489, -1.640043, 0.1895263, 17.29115, 16.96097, 
      3.877544, 4.56585, 5.699979, 13.75763, 13.93032, 5.559056, 5.670705, 
      10.86785, 10.40997, 7.717412, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -1.225706, 11.69911, 
      13.06857, 14.05671, 14.53291, 14.48116, 14.47679, 14.39564, 14.87393, 
      14.7753, 13.68717, 11.97302, 9.113683 ;

   windNorthward = 2.380202, -1.089164, _, -1.794114, 2.936322, _, 2.991843, 
      _, _, 3.023115, _, _, -1.289333, -5.006013, _, -4.117733, _, -7.001625, 
      -8.685597, 3.64881, _, -2.802598, 4.037339, 3.779823, _, -2.583868, 
      3.388475, 2.828758, -2.67919, 2.65556, _, _, -2.773853, _, _, 2.491153, 
      -2.889902, _, -2.150659, _, -14.0447, 0.8029721, _, -12.92819, 
      1.643805, _, 4.388265, 6.986234, 6.684765, 6.673048, -7.191293, 
      -6.860639, 5.680958, 5.309257, 4.528631, -0.4637186, -0.1207601, 
      3.963976, 3.485844, -2.31085, -2.212005, 0.5185826, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      -0.8737034, 1.998885, 1.880142, 1.405234, 0.3026514, -0.5946224, 
      -0.6703909, -2.077407, -5.476562, -6.520739, -11.21046, -12.62324, 
      -9.750257 ;
  } // group GsiHofXBc

group: GsiHofX_linear {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  		string airTemperature:units = "K" ;
  data:

   airTemperature = 217.678, 217.8861, 217.8861, 217.7196, 215.8655, 
      217.1113, 215.7998, 215.6045, 215.8178, 215.8269, 215.8269, 214.962, 
      213.6835, 213.1017, 213.1017, 213.1651, 213.3429, 212.9628, 213.2162, 
      215.9297, 218.5071, 218.4506, 215.8908, 215.8245, 215.8245, 217.3318, 
      215.7757, 215.5481, 216.6158, 215.4153, 215.4153, 216.1747, 216.1477, 
      216.1477, 215.3662, 215.3127, 214.8681, 214.6468, 214.5466, 214.5466, 
      217.6343, 214.7237, 214.9376, 219.8012, 284.4636, _, 285.2984, 
      286.0831, 283.4491, 281.4311, 228.3843, 228.7268, 277.8273, 277.0466, 
      274.6297, 244.1138, 243.209, 271.6857, 269.0067, 254.4606, 255.6868, 
      262.9401, 220.4462, 220.7901, _, 218.8406, 217.6756, 216.2159, 
      211.6913, 212.6143, 229.0036, 227.3472, 213.5354, 212.9029, 211.4324, 
      212.6465, 221.0529, 220.5016, 220.5773, 213.2783, 220.5434, 220.5467, 
      220.5234, 216.0733, 218.9152, _, 218.1147, 218.6232, 218.9254, 
      220.1636, 222.368, 222.8403, 222.9246, 221.1063, 221.0262, 220.6403, 
      219.5535, 218.7283, 212.8596, 212.6263, 213.1989, 214.1484, 215.0985, 
      218.2496, 221.704, 226.1721, 236.6682, 240.4785, 247.9199, 249.9077, 
      257.5207, _, 273.9617, 273.9648, 261.8208, 274.774, 273.1979, 264.5176, 
      267.5702, 219.152, 217.5783, 218.5846, 220.1073, 218.5184, 220.8032, 
      221.8035, 221.8437, 222.2825, 222.715, 228.9698, 230.0241, 227.0518, 
      221.6508, 221.773, 221.7436, 219.4646, 219.5088, 218.348, 213.8849, 
      211.7566, 225.0111, 210.5662, 224.5821, 222.1503, 223.8821, 203.9654, 
      223.6427, 228.243, 208.3333, 202.1172, 203.3788, 211.4454, 225.7168, 
      204.3838, 210.6205, 292.3801, 232.1634, 206.9983, 205.7846, 295.5864, 
      227.5722, 296.1462, 202.0606, 296.2301, 296.2313, 296.2317, 202.6814, 
      201.2967, 236.9904, 236.0444, 237.2904, 200.8362, 244.1877, 232.3323, 
      244.9964, 234.7205, 246.3828, 248.8736, 255.1175, 256.4044, 280.5699, 
      257.1056, 257.2224, 258.2763, 259.7013, 259.8201, 276.4515, 291.1593, 
      221.8936, 226.531, 230.4098, 234.0159, 235.574, 235.7076, 238.2451, 
      244.2239, 244.8024, 247.8318, 249.4795, 252.7007 ;
  } // group GsiHofX_linear

group: GsiQCWeight {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  data:

   airTemperature = _, _, 3.999999, _, _, 3.999999, _, 3.986951, 3.999999, _, 
      3.999999, 3.536047, _, _, 3.999993, _, 3.999999, _, _, _, 3.999999, _, 
      _, _, 3.999999, _, _, _, _, _, 3.999998, 3.999999, _, 3.999999, 
      3.999998, _, _, 3.999997, _, 3.999997, _, _, 3.999998, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3.999998, 3.999998, _, 
      3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999994, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999998, 3.999999, 3.999999, 3.999999, 3.999999, _, 
      3.999999, 3.999998, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999999, 3.999999, 3.999999, 3.999999, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3.999999, 3.999999, 3.999998, 
      3.999999, 3.999999, 3.999999, 3.999722, 3.999688, 3.999879, 3.999999, 
      3.999993, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 3.999526, 3.99914, 3.998858, 3.998767, 
      3.998995, 3.999021, 3.999238, 3.999388, 3.999463, 3.999646, 3.999655, 
      3.999672, 3.999651, _, 3.998883, 3.998775, 3.99964, 3.999556, 3.99958, 
      3.999678, 3.999619, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, 3.999686, 3.99967, 3.999628, 3.999677, 3.99959, 3.999672, 3.999681, 
      3.999685, 3.999655, 3.999685, 3.999668, 3.999559, 3.999662, 3.99966, 
      3.999681, 3.999686, 3.999635, 3.999674, 3.999686, 3.999568, 3.999585, 
      3.999605, 3.999686, 3.999686, 3.999686, 3.999677, 3.999685, 3.999686, 
      3.999686, 3.999675, 3.999675, 3.999685, 3.999686, 3.998787, 3.999668, 
      3.99968, 3.999686, 3.999686, 3.999686, 3.999686, 3.999681, 3.997346, 
      3.992576, 3.999686, 3.998926, 3.999177, 3.99968, 3.999667, 3.99966, 
      3.999683, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 3.999565, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      3.999598, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      3.999274, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 3.999591, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 3.999999, 3.999999, _, 3.999998, 3.999931, _, 3.999999, _, 
      _, 3.999999, _, _, 3.999998, 3.999998, _, 3.999994, _, 3.999995, 
      3.999998, 3.999987, _, 3.999999, 3.999945, 3.999999, _, 3.998322, 
      3.999998, 3.999992, 3.999999, 3.999996, _, _, 3.999999, _, _, 3.999434, 
      3.999997, _, 3.999999, _, 3.999972, 3.999991, _, 3.999999, 3.999999, _, 
      3.999999, 3.999992, 3.999884, 3.999978, 3.999998, 3.999998, 3.999996, 
      3.999997, 3.999999, 3.999999, 3.999999, 3.999985, 3.999998, 3.999998, 
      3.999999, 3.999999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999998, 3.999996 ;

   windNorthward = 3.999999, 3.999999, _, 3.999998, 3.999931, _, 3.999999, _, 
      _, 3.999999, _, _, 3.999998, 3.999998, _, 3.999994, _, 3.999995, 
      3.999998, 3.999987, _, 3.999999, 3.999945, 3.999999, _, 3.998322, 
      3.999998, 3.999992, 3.999999, 3.999996, _, _, 3.999999, _, _, 3.999434, 
      3.999997, _, 3.999999, _, 3.999972, 3.999991, _, 3.999999, 3.999999, _, 
      3.999999, 3.999992, 3.999884, 3.999978, 3.999998, 3.999998, 3.999996, 
      3.999997, 3.999999, 3.999999, 3.999999, 3.999985, 3.999998, 3.999998, 
      3.999999, 3.999999, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 3.999999, 
      3.999999, 3.999998, 3.999996 ;
  } // group GsiQCWeight

group: GsiUseFlag {
  variables:
  	int airTemperature(Location) ;
  		airTemperature:_FillValue = -2147483647 ;
  	int specificHumidity(Location) ;
  		specificHumidity:_FillValue = -2147483647 ;
  	int stationPressure(Location) ;
  		stationPressure:_FillValue = -2147483647 ;
  	int windEastward(Location) ;
  		windEastward:_FillValue = -2147483647 ;
  	int windNorthward(Location) ;
  		windNorthward:_FillValue = -2147483647 ;
  data:

   airTemperature = _, _, 1, _, _, 1, _, 1, 1, _, 1, 1, _, _, 1, _, 1, _, _, 
      _, 1, _, _, _, 1, _, _, _, _, _, 1, 1, _, 1, 1, _, _, 1, _, 1, _, _, 1, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, 1, _, 1, 1, 
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, 1, 1, 1, 1, 1, 
      1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, -1, -1, -1, -1, -1, -1, -1, -1, 1, 1, 1, 1, 1, 
      _, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
      -1, -1, 1, -1, -1, -1, 1, -1, 1, -1, 1, 1, 1, -1, -1, -1, -1, -1, -1, 
      -1, -1, 1, -1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 
      _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 1, 1, _, 1, 1, _, 1, _, _, 1, _, _, 1, 1, _, 1, _, 1, 1, 1, 
      _, 1, 1, 1, _, 1, 1, 1, 1, 1, _, _, 1, _, _, 1, 1, _, 1, _, 1, 1, _, 1, 
      1, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, 
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

   windNorthward = 1, 1, _, 1, 1, _, 1, _, _, 1, _, _, 1, 1, _, 1, _, 1, 1, 
      1, _, 1, 1, 1, _, 1, 1, 1, 1, 1, _, _, 1, _, _, 1, 1, _, 1, _, 1, 1, _, 
      1, 1, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;
  } // group GsiUseFlag

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -2208988800LL ;
  		string dateTime:units = "seconds since 1970-01-01T00:00:00Z" ;
  	float height(Location) ;
  		height:_FillValue = 9.96921e+36f ;
  		string height:units = "m" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  		string latitude:units = "degrees_north" ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  		string longitude:units = "degrees_east" ;
  	float pressure(Location) ;
  		pressure:_FillValue = 9.96921e+36f ;
  		string pressure:units = "Pa" ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  	float stationElevation(Location) ;
  		stationElevation:_FillValue = 9.96921e+36f ;
  		string stationElevation:units = "m" ;
  	string stationIdentification(Location) ;
  		string stationIdentification:_FillValue = "" ;
  data:

   dateTime = 1523750874, 1523750682, 1523750682, 1523750656, 1523751089, 
      1523750615, 1523751161, 1523750559, 1523751185, 1523751198, 1523751198, 
      1523750536, 1523750491, 1523750395, 1523750395, 1523750415, 1523750470, 
      1523750350, 1523750318, 1523751353, 1523753617, 1523753609, 1523751540, 
      1523751650, 1523751650, 1523753440, 1523751756, 1523751996, 1523753319, 
      1523752078, 1523752078, 1523753240, 1523753234, 1523753234, 1523752109, 
      1523752138, 1523752882, 1523752772, 1523752720, 1523752720, 1523750105, 
      1523752394, 1523752316, 1523750036, 1523747951, 1523747951, 1523747971, 
      1523748008, 1523748102, 1523748153, 1523749796, 1523749787, 1523748241, 
      1523748262, 1523748340, 1523749374, 1523749398, 1523748450, 1523748553, 
      1523749105, 1523749072, 1523748794, 1523753931, 1523747807, 1523747807, 
      1523747807, 1523747807, 1523747807, 1523747807, 1523747807, 1523747807, 
      1523747807, 1523747807, 1523753053, 1523752551, 1523751915, 1523749704, 
      1523749873, 1523749942, 1523751495, 1523750129, 1523750161, 1523750187, 
      1523751049, 1523750531, 1523748600, 1523750710, 1523750787, 1523750828, 
      1523750930, 1523751114, 1523751209, 1523751490, 1523751990, 1523752016, 
      1523752474, 1523752910, 1523753312, 1523750637, 1523750542, 1523750464, 
      1523750424, 1523750386, 1523750288, 1523750194, 1523750082, 1523749808, 
      1523749702, 1523749492, 1523749439, 1523749238, 1523748528, 1523748528, 
      1523748546, 1523749101, 1523748629, 1523748681, 1523748986, 1523748832, 
      1523752198, 1523753031, 1523752628, 1523751740, 1523753284, 1523753654, 
      1523753804, 1523753810, 1523753896, 1523753997, 1523754909, 1523755022, 
      1523754710, 1523751214, 1523750840, 1523750835, 1523750552, 1523750405, 
      1523755503, 1523755182, 1523755053, 1523756170, 1523754978, 1523756126, 
      1523755875, 1523756058, 1523753797, 1523756031, 1523756503, 1523754865, 
      1523753918, 1523754606, 1523753534, 1523753191, 1523754686, 1523753557, 
      1523751049, 1523756955, 1523754813, 1523754767, 1523750931, 1523753126, 
      1523750902, 1523754341, 1523750880, 1523750871, 1523750867, 1523754465, 
      1523754231, 1523752578, 1523752641, 1523757525, 1523754043, 1523752305, 
      1523752891, 1523752279, 1523752736, 1523752235, 1523752157, 1523751960, 
      1523751926, 1523751375, 1523751908, 1523751905, 1523751878, 1523751843, 
      1523751840, 1523751471, 1523749372, 1523750501, 1523750501, 1523750501, 
      1523750501, 1523750501, 1523750501, 1523750501, 1523750501, 1523750501, 
      1523750501, 1523750501, 1523750501 ;

   height = 0, 0, 13700, 0, 0, _, 0, _, _, 0, 16280, _, 0, 0, _, 0, _, 0, 0, 
      0, _, 0, 0, 0, 18540, 0, 0, 0, 0, 0, 20680, _, 0, 26460, _, 0, 0, _, 0, 
      23890, 0, 0, _, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 30620, _, 2, _, _, _, _, _, _, _, _, 26230, 23720, 20540, _, 10330, 
      _, 18440, _, 11770, _, 16210, 13620, 100, _, _, 9910, _, 11340, _, 
      13220, _, 15850, 18140, 20320, _, _, _, _, 10160, _, _, 9010, _, 7080, 
      _, 5500, _, _, 675, 675, 765, _, _, 1443, 2968, _, 18220, _, 20370, 
      15930, 23650, _, 26250, _, _, _, _, _, 30780, 13300, 11430, _, 9990, _, 
      23790, _, _, _, _, _, _, _, _, 26430, _, 20600, _, _, _, 12230, _, 
      14060, 1518, 31050, _, _, _, _, 786, _, _, _, 612, 18600, _, _, 9480, 
      33900, 16490, _, 10730, _, _, 7450, _, _, _, 3149, _, 5800, _, _, _, _, 
      6286.768, 6286.768, 6286.768, 6286.768, 6286.768, 6286.768, 6286.768, 
      6286.768, 6286.768, 6286.768, 6286.768, 6286.768, 6286.768 ;

   latitude = 44.77628, 44.77816, 44.77816, 44.77919, 44.78084, 44.78087, 
      44.78238, 44.78266, 44.78277, 44.78301, 44.78301, 44.78324, 44.78408, 
      44.78418, 44.78418, 44.78419, 44.78431, 44.7851, 44.78624, 44.78827, 
      44.79156, 44.79156, 44.79337, 44.79533, 44.79533, 44.7964, 44.79758, 
      44.79822, 44.79937, 44.80019, 44.80019, 44.80055, 44.80065, 44.80065, 
      44.80207, 44.80409, 44.80432, 44.80521, 44.80585, 44.80585, 44.81009, 
      44.81119, 44.81156, 44.82153, 44.83, 44.83, 44.83075, 44.83342, 
      44.84194, 44.84638, 44.84642, 44.8469, 44.85229, 44.85331, 44.85671, 
      44.85708, 44.85708, 44.86032, 44.86301, 44.86345, 44.86498, 44.86869, 
      54.73114, 54.75, 54.75, 54.75, 54.75, 54.75, 54.75, 54.75, 54.75, 
      54.75, 54.75, 54.80032, 54.8373, 54.87028, 54.87428, 54.88316, 
      54.88366, 54.88514, 54.89388, 54.89465, 54.89529, 54.90061, 54.90599, 
      62.08, 68.69463, 68.69873, 68.70068, 68.70525, 68.71354, 68.71751, 
      68.73039, 68.75166, 68.75278, 68.77066, 68.79052, 68.80064, 50.15633, 
      50.17497, 50.19108, 50.19964, 50.20792, 50.2281, 50.24597, 50.26628, 
      50.31132, 50.32695, 50.35397, 50.35933, 50.37483, 50.38, 50.38, 
      50.38016, 50.38275, 50.38363, 50.38607, 50.38754, 50.39029, 53.48677, 
      53.48981, 53.49107, 53.49156, 53.49279, 53.50296, 53.50717, 53.50733, 
      53.50936, 53.51147, 53.51159, 53.51183, 53.51622, 53.5168, 53.55087, 
      53.55141, 53.58424, 53.60339, 24.90497, 24.90725, 24.91282, 24.91628, 
      24.91748, 24.91795, 24.91933, 24.9194, 24.9195, 24.9199, 24.92107, 
      24.92585, 24.92602, 24.92676, 24.92727, 24.92738, 24.92807, 24.92822, 
      24.92888, 24.92899, 24.92925, 24.92954, 24.9297, 24.92986, 24.92993, 
      24.92994, 24.92999, 24.93, 24.93, 24.9309, 24.93496, 24.93516, 
      24.93546, 24.9367, 24.93723, 24.93774, 24.93776, 24.93785, 24.93801, 
      24.93897, 24.94201, 24.94674, 24.94722, 24.94744, 24.94775, 24.94786, 
      24.94907, 24.95046, 24.95055, 24.9531, 16.9616, 16.96161, 16.96161, 
      16.96161, 16.96161, 16.96161, 16.96161, 16.96161, 16.96161, 16.96161, 
      16.96161, 16.96161, 16.96161 ;

   longitude = 359.7401, 359.7238, 359.7238, 359.7203, 359.7608, 359.7143, 
      359.7675, 359.7045, 359.7682, 359.7686, 359.7686, 359.6998, 359.6899, 
      359.6703, 359.6703, 359.6738, 359.6851, 359.6638, 359.6594, 359.7689, 
      359.894, 359.894, 359.7762, 359.7842, 359.7842, 359.8686, 359.7866, 
      359.7947, 359.853, 359.7992, 359.7992, 359.8475, 359.8472, 359.8472, 
      359.7999, 359.7994, 359.8347, 359.8323, 359.8304, 359.8304, 359.5946, 
      359.8074, 359.8012, 359.5667, 359.32, 359.32, 359.3195, 359.318, 
      359.3169, 359.3186, 359.5021, 359.5006, 359.3242, 359.326, 359.3319, 
      359.4338, 359.4377, 359.3364, 359.3397, 359.3927, 359.3881, 359.3561, 
      18.21814, 17.53, 17.53, 17.53, 17.53, 17.53, 17.53, 17.53, 17.53, 
      17.53, 17.53, 18.17319, 18.15634, 18.11426, 17.91357, 17.95114, 
      17.95688, 18.08035, 17.97266, 17.97495, 17.97623, 18.04828, 18.00333, 
      129.75, 160.6873, 160.6581, 160.6475, 160.6257, 160.5861, 160.5676, 
      160.537, 160.503, 160.5021, 160.4753, 160.443, 160.4069, 116.6575, 
      116.6497, 116.643, 116.6394, 116.6359, 116.6263, 116.6168, 116.6066, 
      116.5862, 116.5797, 116.5671, 116.5652, 116.5527, 116.52, 116.52, 
      116.5195, 116.5492, 116.5237, 116.5287, 116.5473, 116.5389, 127.3618, 
      127.4372, 127.4029, 127.309, 127.4524, 127.464, 127.4667, 127.4668, 
      127.4687, 127.4714, 127.5126, 127.5137, 127.5078, 127.2558, 127.2378, 
      127.2376, 127.2306, 127.2292, 47.6329, 47.63748, 47.64288, 47.63132, 
      47.64453, 47.62943, 47.62592, 47.6261, 47.47165, 47.62573, 47.64197, 
      47.64374, 47.51379, 47.633, 47.34253, 47.16083, 47.63541, 47.35529, 
      46.71042, 47.65985, 47.64236, 47.64023, 46.71722, 47.12946, 46.71909, 
      47.61295, 46.71988, 46.72, 46.72, 47.62079, 47.59763, 46.91943, 46.935, 
      47.63739, 47.5549, 46.86407, 47.03003, 46.85919, 46.96704, 46.85165, 
      46.83902, 46.81018, 46.8056, 46.7218, 46.80292, 46.80246, 46.79858, 
      46.79312, 46.79263, 46.73419, 73.33868, 73.33868, 73.33868, 73.33868, 
      73.33868, 73.33868, 73.33868, 73.33868, 73.33868, 73.33868, 73.33868, 
      73.33868, 73.33868 ;

   pressure = 12900, 15000, 15000, 15300, 10900, 15800, 10300, 16500, 10100, 
      10000, 10000, 16800, 17400, 18800, 18800, 18500, 17700, 19500, 20000, 
      8850, 1480, 1490, 7640, 7000, 7000, 1700, 6440, 5330, 1870, 5000, 5000, 
      1990, 2000, 2000, 4880, 4770, 2640, 2880, 3000, 3000, 23700, 3890, 
      4140, 25000, 101100, 101100, 100000, 97800, 92500, 89700, 30000, 30200, 
      85000, 83900, 80000, 40700, 40000, 74700, 70000, 48900, 50000, 60000, 
      1000, 1000, 101900, 1150, 1270, 1440, 2470, 4650, 650, 700, 7240, 2000, 
      3000, 5000, 28500, 25000, 23700, 7000, 20500, 20000, 19600, 10000, 
      15000, 99600, 27400, 25800, 25000, 23100, 20000, 18600, 15000, 10200, 
      10000, 7000, 5000, 3660, 21000, 22700, 24200, 25000, 25800, 27900, 
      30000, 32700, 40000, 43200, 50000, 51900, 59400, 93600, 93600, 92500, 
      65000, 87800, 85000, 70000, 77300, 7000, 3650, 5000, 10000, 3000, 2250, 
      2000, 1990, 1860, 1720, 860, 790, 1000, 15000, 20000, 20100, 25000, 
      28000, 3000, 3870, 4290, 1800, 4560, 1860, 2250, 1960, 12300, 2000, 
      1400, 5000, 11100, 6210, 15300, 20000, 5800, 15000, 85000, 1000, 5220, 
      5420, 91000, 21000, 92500, 7770, 93400, 93900, 94100, 7000, 8520, 
      31400, 30000, 660, 10000, 38100, 25000, 38800, 28000, 40000, 42200, 
      48200, 49300, 70000, 49900, 50000, 50900, 52100, 52200, 66000, 78900, 
      20270, 22000, 23510, 25000, 25700, 25760, 26900, 30000, 30550, 33600, 
      35600, 38250 ;

   sequenceNumber = 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 
      29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 
      29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 
      29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 53, 53, 53, 53, 53, 53, 
      53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 
      115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 65, 
      65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 160, 65, 65, 65, 65, 
      65, 65, 65, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 
      160, 160, 160, 160, 160, 160, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 
      91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 
      91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 
      91, 91, 91, 91, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 
      255, 255 ;

   stationElevation = 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
      47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
      47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
      47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 2, 2, 2, 2, 2, 2, 2, 2, 
      2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 100, 26, 26, 26, 26, 26, 
      26, 26, 26, 26, 26, 26, 26, 675, 675, 675, 675, 675, 675, 675, 675, 
      675, 675, 675, 675, 675, 675, 675, 675, 675, 675, 675, 675, 675, 228, 
      228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 228, 
      228, 228, 228, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 
      612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 
      612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 
      612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 612, 34, 34, 34, 34, 
      34, 34, 34, 34, 34, 34, 34, 34, 34 ;

   stationIdentification = "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "07510", "07510", "07510", "07510", "07510", "07510", "07510", 
      "07510", "12120", "12120", "12120", "12120", "12120", "12120", "12120", 
      "12120", "12120", "12120", "12120", "12120", "12120", "12120", "12120", 
      "12120", "12120", "12120", "12120", "12120", "12120", "12120", "12120", 
      "24959", "25123", "25123", "25123", "25123", "25123", "25123", "25123", 
      "25123", "25123", "25123", "25123", "25123", "30965", "30965", "30965", 
      "30965", "30965", "30965", "30965", "30965", "30965", "30965", "30965", 
      "30965", "30965", "30965", "30965", "30965", "30965", "30965", "30965", 
      "30965", "30965", "31300", "31300", "31300", "31300", "31300", "31300", 
      "31300", "31300", "31300", "31300", "31300", "31300", "31300", "31300", 
      "31300", "31300", "31300", "31300", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "40437", "40437", 
      "40437", "40437", "40437", "40437", "40437", "40437", "43110", "43110", 
      "43110", "43110", "43110", "43110", "43110", "43110", "43110", "43110", 
      "43110", "43110", "43110" ;
  } // group MetaData

group: ObsError {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  		string airTemperature:units = "K" ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  		string specificHumidity:units = "1" ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  		string stationPressure:units = "Pa" ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  		string windEastward:units = "m s-1" ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  		string windNorthward:units = "m s-1" ;
  data:

   airTemperature = _, _, 1, _, _, 1, _, 1.1, 0.8, _, 0.8, 1.1, _, _, 1.2, _, 
      1.1, _, _, _, 1.4, _, _, _, 0.8, _, _, _, _, _, 0.9, 1.3, _, 1.3, 0.9, 
      _, _, 1, _, 1, _, _, 0.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, 1.5, 1.5, _, 1.5, 1.4, 1.4, 1.1, 0.9, 1.5, 1.5, 0.8, 1.3, 
      1, 0.9, 1, 1.2, 1.2, 0.8, 1.2, 1.2, 1.2, 0.8, 1, _, 1.1, 1.2, 1.2, 1.2, 
      1.2, 1.1, 1, 0.8, 0.8, 0.8, 0.9, 1, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, 0.8, 1, 0.9, 0.8, 1, 1.2, 1.3, 1.3, 1.3, 
      1.3, 1.5, 1.5, 1.5, 1, 1.2, 1.2, 1.2, 1, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 1.056813e-05, 9.957423e-06, 1.009526e-05, 
      1.106756e-05, 1.200879e-05, 1.653376e-05, 2.317654e-05, 3.509987e-05, 
      8.544992e-05, 0.0001147122, 0.0001975877, 0.0002286237, 0.0003814484, 
      _, 0.0008766068, 0.0008767928, 0.0004945507, 0.0009753293, 
      0.0008994794, 0.0005680757, 0.0006505361, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 1.431543e-05, 1.110419e-05, 1.003266e-05, 
      2.407659e-05, 9.466662e-06, 2.328926e-05, 1.919881e-05, 2.204181e-05, 
      5.867995e-06, 2.162867e-05, 3.104534e-05, 8.654431e-06, 5.022742e-06, 
      6.947986e-06, 1.2853e-05, 5.41556e-05, 7.45339e-06, 1.196863e-05, 
      0.003287753, 4.396388e-05, 8.303241e-06, 7.985352e-06, 0.0037453, 
      6.315239e-05, 0.003812299, 5.541402e-06, 0.003801987, 0.003802242, 
      0.003802343, 6.162792e-06, 5.046217e-06, 0.0001117017, 0.0001065203, 
      6.678051e-05, 4.642167e-06, 0.0001840855, 8.748625e-05, 0.0001960853, 
      9.978229e-05, 0.0002161481, 0.0002566602, 0.0003862471, 0.0004218426, 
      0.001844437, 0.0004408921, 0.0004440425, 0.0004738013, 0.0005239225, 
      0.0005280467, 0.001465403, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 2.3, 2.4, _, 2.4, 2.2, _, 2.1, _, _, 2.1, _, _, 2.5, 2.6, 
      _, 2.6, _, 2.7, 2.7, 2.1, _, 2.1, 2.1, 2.1, _, 2.1, 2.1, 2.1, 2.1, 2.1, 
      _, _, 2.1, _, _, 2.1, 2.1, _, 2.1, _, 3.1, 2.1, _, 3.2, 1.4, _, 1.4, 
      1.4, 1.5, 1.5, 3, 3, 1.5, 1.5, 1.6, 2.6, 2.6, 1.6, 1.6, 2.1, 2.1, 1.9, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 1.6, 2.7, 2.9, 3.1, 3.2, 3.2, 3.2, 3.1, 3, 3, 2.9, 2.8, 
      2.7 ;

   windNorthward = 2.3, 2.4, _, 2.4, 2.2, _, 2.1, _, _, 2.1, _, _, 2.5, 2.6, 
      _, 2.6, _, 2.7, 2.7, 2.1, _, 2.1, 2.1, 2.1, _, 2.1, 2.1, 2.1, 2.1, 2.1, 
      _, _, 2.1, _, _, 2.1, 2.1, _, 2.1, _, 3.1, 2.1, _, 3.2, 1.4, _, 1.4, 
      1.4, 1.5, 1.5, 3, 3, 1.5, 1.5, 1.6, 2.6, 2.6, 1.6, 1.6, 2.1, 2.1, 1.9, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 1.6, 2.7, 2.9, 3.1, 3.2, 3.2, 3.2, 3.1, 3, 3, 2.9, 2.8, 
      2.7 ;
  } // group ObsError

group: ObsType {
  variables:
  	int airTemperature(Location) ;
  		airTemperature:_FillValue = -2147483647 ;
  	int specificHumidity(Location) ;
  		specificHumidity:_FillValue = -2147483647 ;
  	int stationPressure(Location) ;
  		stationPressure:_FillValue = -2147483647 ;
  	int windEastward(Location) ;
  		windEastward:_FillValue = -2147483647 ;
  	int windNorthward(Location) ;
  		windNorthward:_FillValue = -2147483647 ;
  data:

   airTemperature = _, _, 120, _, _, 120, _, 120, 120, _, 120, 120, _, _, 
      120, _, 120, _, _, _, 120, _, _, _, 120, _, _, _, _, _, 120, 120, _, 
      120, 120, _, _, 120, _, 120, _, _, 120, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, 120, 120, _, 120, 120, 120, 120, 120, 120, 
      120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      _, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 120, 120, 120, 
      120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      120, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      120, 120, 120, 120, _, 120, 120, 120, 120, 120, 120, 120, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, 120, 120, 120, 120, 120, 120, 
      120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 
      120, 120, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 120, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 120, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 120, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      120, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 220, 220, _, 220, 220, _, 220, _, _, 220, _, _, 220, 220, 
      _, 220, _, 220, 220, 220, _, 220, 220, 220, _, 220, 220, 220, 220, 220, 
      _, _, 220, _, _, 220, 220, _, 220, _, 220, 220, _, 220, 220, _, 220, 
      220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 
      220, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 
      220, 220, 220 ;

   windNorthward = 220, 220, _, 220, 220, _, 220, _, _, 220, _, _, 220, 220, 
      _, 220, _, 220, 220, 220, _, 220, 220, 220, _, 220, 220, 220, 220, 220, 
      _, _, 220, _, _, 220, 220, _, 220, _, 220, 220, _, 220, 220, _, 220, 
      220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 
      220, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 
      220, 220, 220 ;
  } // group ObsType

group: ObsValue {
  variables:
  	float airTemperature(Location) ;
  		airTemperature:_FillValue = 9.96921e+36f ;
  		string airTemperature:units = "K" ;
  	float specificHumidity(Location) ;
  		specificHumidity:_FillValue = 9.96921e+36f ;
  		string specificHumidity:units = "1" ;
  	float stationPressure(Location) ;
  		stationPressure:_FillValue = 9.96921e+36f ;
  		string stationPressure:units = "Pa" ;
  	float windEastward(Location) ;
  		windEastward:_FillValue = 9.96921e+36f ;
  		string windEastward:units = "m s-1" ;
  	float windNorthward(Location) ;
  		windNorthward:_FillValue = 9.96921e+36f ;
  		string windNorthward:units = "m s-1" ;
  data:

   airTemperature = _, _, 217.85, _, _, 217.85, _, 220.45, 216.65, _, 216.65, 
      220.65, _, _, 210.45, _, 213.05, _, _, _, 219.05, _, _, _, 216.65, _, 
      _, _, _, _, 216.65, 215.45, _, 215.45, 216.65, _, _, 216.45, _, 216.25, 
      _, _, 213.45, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      218.25, 218.25, _, 219.85, 216.05, 217.45, 210.45, 213.45, 228.45, 
      228.85, 211.85, 212.85, 211.85, 212.45, 220.65, 220.05, 219.25, 212.45, 
      222.45, 221.05, 220.05, 216.45, 218.65, _, 216.65, 220.25, 220.25, 
      218.65, 222.25, 223.05, 221.65, 220.85, 221.25, 220.45, 220.05, 219.05, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 219.85, 
      217.45, 219.85, 219.85, 219.25, 220.45, 217.25, 217.25, 218.05, 222.45, 
      225.65, 228.45, 225.05, 221.85, 222.05, 222.05, 220.65, 218.65, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 3e-06, 2e-06, 3e-06, 3e-06, 5e-06, 7e-06, 
      1.4e-05, 2.8e-05, 8.5e-05, 0.000175, 0.000227, 0.000238, 0.000106, _, 
      0.000896, 0.000846, 0.000238, 0.000997, 0.000881, 0.000619, 0.00075, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3e-06, 2e-06, 1e-06, 
      1.1e-05, 1e-06, 1.2e-05, 8e-06, 7e-06, 1e-06, 7e-06, 1.6e-05, 1e-06, 
      1e-06, 1e-06, 2e-06, 2e-06, 1e-06, 1e-06, 0.004482, 4.2e-05, 1e-06, 
      1e-06, 0.004372, 3e-06, 0.004557, 1e-06, 0.004713, 0.004893, 0.004745, 
      1e-06, 1e-06, 9e-06, 1.1e-05, 0.000117, 1e-06, 1.9e-05, 5e-06, 7.4e-05, 
      7e-06, 9.6e-05, 0.000112, 0.00029, 0.000377, 0.003583, 0.000935, 
      0.001041, 0.001826, 0.002373, 0.002428, 0.00306, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 101100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      101900, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      99600, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, 93600, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 3.3, 10.1, _, 10.7, 12, _, 2.7, _, _, 2.2, _, _, 18.4, 
      13.3, _, 14.8, _, 9.2, 13.1, -1.9, _, 9.5, 8.2, 3.3, _, 14.4, 0.3, 5, 
      6, 3.6, _, _, 4.8, _, _, -3, 0.8, _, 3.3, _, 34.8, 7.9, _, 29.4, -1.8, 
      _, -2.6, -3.7, 1.8, 3.3, 13, 12.6, 6.7, 7.2, 4.7, 12.9, 12.9, 1.8, 3.3, 
      11.2, 10.7, 7.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, 0.3, 10.4, 12.1, 13.3, 14.4, 14.4, 
      14.9, 14.5, 13, 13.9, 14.7, 13.6, 10.3 ;

   windNorthward = 1.5, -3.7, _, -5, 3.2, _, 1.5, _, _, 2.2, _, _, -1.6, 
      -1.2, _, 1.3, _, -3.3, -4.8, 5.4, _, -2.5, 0.7, 3.3, _, -3.9, 1.5, 
      -0.9, -1.6, 6.2, _, _, -1.7, _, _, 8.3, -0.6, _, -1.5, _, -20.1, -2.1, 
      _, -17, 3.1, _, 5.6, 10.1, 10.1, 9.2, -6.1, -5.9, 5.7, 5, 4.7, 0, 0, 
      2.5, 3.3, -5.2, -5, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, 0.3, 2.8, 4.4, 1.2, 0, 0, 0, 
      -5.3, -6.1, -8, -8.5, -16.2, -14.7 ;
  } // group ObsValue

group: PreQC {
  variables:
  	int airTemperature(Location) ;
  		airTemperature:_FillValue = -2147483647 ;
  	int specificHumidity(Location) ;
  		specificHumidity:_FillValue = -2147483647 ;
  	int stationPressure(Location) ;
  		stationPressure:_FillValue = -2147483647 ;
  	int windEastward(Location) ;
  		windEastward:_FillValue = -2147483647 ;
  	int windNorthward(Location) ;
  		windNorthward:_FillValue = -2147483647 ;
  data:

   airTemperature = _, _, 2, _, _, 2, _, 2, 2, _, 2, 2, _, _, 2, _, 2, _, _, 
      _, 2, _, _, _, 2, _, _, _, _, _, 2, 2, _, 2, 2, _, _, 2, _, 2, _, _, 2, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, _, 2, 2, 
      2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, 2, 
      2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 9, 9, 9, 9, 9, 9, 15, 15, 2, 2, 2, 2, 2, _, 2, 
      2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 2, 9, 9, 9, 2, 9, 
      2, 9, 2, 2, 2, 9, 9, 15, 15, 9, 9, 15, 9, 2, 9, 2, 2, 2, 2, 2, 2, 2, 2, 
      2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 2, 2, _, 2, 2, _, 2, _, _, 2, _, _, 2, 2, _, 2, _, 2, 2, 2, 
      _, 2, 2, 2, _, 2, 2, 2, 2, 2, _, _, 2, _, _, 2, 2, _, 2, _, 2, 2, _, 2, 
      2, _, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 
      2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

   windNorthward = 2, 2, _, 2, 2, _, 2, _, _, 2, _, _, 2, 2, _, 2, _, 2, 2, 
      2, _, 2, 2, 2, _, 2, 2, 2, 2, 2, _, _, 2, _, _, 2, 2, _, 2, _, 2, 2, _, 
      2, 2, _, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;
  } // group PreQC

group: PreUseFlag {
  variables:
  	int airTemperature(Location) ;
  		airTemperature:_FillValue = -2147483647 ;
  	int specificHumidity(Location) ;
  		specificHumidity:_FillValue = -2147483647 ;
  	int stationPressure(Location) ;
  		stationPressure:_FillValue = -2147483647 ;
  	int windEastward(Location) ;
  		windEastward:_FillValue = -2147483647 ;
  	int windNorthward(Location) ;
  		windNorthward:_FillValue = -2147483647 ;
  data:

   airTemperature = _, _, 0, _, _, 0, _, 0, 0, _, 0, 0, _, _, 0, _, 0, _, _, 
      _, 0, _, _, _, 0, _, _, _, _, _, 0, 0, _, 0, 0, _, _, 0, _, 0, _, _, 0, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   specificHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, 101, 101, 101, 101, 101, 101, 101, 101, 0, 0, 
      0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 
      101, 101, 101, 101, 101, 101, 101, 0, 101, 101, 101, 0, 101, 0, 101, 0, 
      0, 0, 101, 101, 101, 101, 101, 101, 101, 101, 0, 101, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   stationPressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _ ;

   windEastward = 0, 0, _, 0, 0, _, 0, _, _, 0, _, _, 0, 0, _, 0, _, 0, 0, 0, 
      _, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, 0, _, _, 0, 0, _, 0, _, 0, 0, _, 0, 
      0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

   windNorthward = 0, 0, _, 0, 0, _, 0, _, _, 0, _, _, 0, 0, _, 0, _, 0, 0, 
      0, _, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, 0, _, _, 0, 0, _, 0, _, 0, 0, _, 
      0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreUseFlag
}
