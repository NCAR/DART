netcdf sgpswatsE13.b1 {
dimensions:
	time = UNLIMITED ; // (1824 currently)
	depth = 8 ;
variables:
	int base_time ;
		base_time:string = "1-May-2003,0:07:00 GMT" ;
		base_time:long_name = "Base time in Epoch" ;
		base_time:units = "seconds since 1970-1-1 0:00:00 0:00" ;
	double time_offset(time) ;
		time_offset:long_name = "Time offset from base_time" ;
		time_offset:units = "seconds since 2003-05-01 00:07:00 0:00" ;
	int depth(depth) ;
		depth:long_name = "Sensor Depth below surface" ;
		depth:units = "cm" ;
	float tref(time) ;
		tref:long_name = "Reference Thermistor Temperature" ;
		tref:units = "degC" ;
		tref:valid_min = -25.f ;
		tref:valid_max = 50.f ;
		tref:valid_delta = 20.f ;
		tref:resolution = 0.1f ;
		tref:missing_value = -9999.f ;
		tref:accuracy = "0.2 degC" ;
	int qc_tref(time) ;
		qc_tref:long_name = "Quality check results on field: Reference Thermistor Temperature" ;
		qc_tref:units = "unitless" ;
	float tsoil_W(time, depth) ;
		tsoil_W:long_name = "Soil Temperature, West Profile" ;
		tsoil_W:units = "degC" ;
		tsoil_W:valid_min = -20.f ;
		tsoil_W:valid_max = 50.f ;
		tsoil_W:valid_delta = 20.f ;
		tsoil_W:resolution = 0.1f ;
		tsoil_W:missing_value = -9999.f ;
		tsoil_W:accuracy = "0.5 degC" ;
	int qc_tsoil_W(time, depth) ;
		qc_tsoil_W:long_name = "Quality check results on field: Soil Temperature, West Profile" ;
		qc_tsoil_W:units = "unitless" ;
	float trise_W(time, depth) ;
		trise_W:long_name = "Sensor Temperature Rise, West Profile" ;
		trise_W:units = "degC" ;
		trise_W:valid_min = 1.f ;
		trise_W:valid_max = 4.5f ;
		trise_W:valid_delta = 3.5f ;
		trise_W:resolution = 0.01f ;
		trise_W:missing_value = -9999.f ;
		trise_W:accuracy = "0.04 degC" ;
	int qc_trise_W(time, depth) ;
		qc_trise_W:long_name = "Quality check results on field: Sensor Temperature Rise, West Profile" ;
		qc_trise_W:units = "unitless" ;
	float soilwatpot_W(time, depth) ;
		soilwatpot_W:long_name = "Soil Water Potential, West Profile" ;
		soilwatpot_W:units = "kPa" ;
		soilwatpot_W:valid_min = -7000.f ;
		soilwatpot_W:valid_max = 0.f ;
		soilwatpot_W:valid_delta = 7000.f ;
		soilwatpot_W:missing_value = -9999.f ;
	int qc_soilwatpot_W(time, depth) ;
		qc_soilwatpot_W:long_name = "Quality check results on field: Soil Water Potential, West Profile" ;
		qc_soilwatpot_W:units = "unitless" ;
	float watcont_W(time, depth) ;
		watcont_W:long_name = "Volumetric Water Content, West Profile" ;
		watcont_W:units = "m3/m3" ;
		watcont_W:valid_min = 0.f ;
		watcont_W:valid_max = 0.55f ;
		watcont_W:valid_delta = 0.55f ;
		watcont_W:missing_value = -9999.f ;
	int qc_watcont_W(time, depth) ;
		qc_watcont_W:long_name = "Quality check results on field: Volumetric Water Content, West Profile" ;
		qc_watcont_W:units = "unitless" ;
	float tsoil_E(time, depth) ;
		tsoil_E:long_name = "Soil Temperature, East Profile" ;
		tsoil_E:units = "degC" ;
		tsoil_E:valid_min = -20.f ;
		tsoil_E:valid_max = 50.f ;
		tsoil_E:valid_delta = 20.f ;
		tsoil_E:resolution = 0.1f ;
		tsoil_E:missing_value = -9999.f ;
		tsoil_E:accuracy = "0.5 degC" ;
	int qc_tsoil_E(time, depth) ;
		qc_tsoil_E:long_name = "Quality check results on field: Soil Temperature, East Profile" ;
		qc_tsoil_E:units = "unitless" ;
	float trise_E(time, depth) ;
		trise_E:long_name = "Sensor Temperature Rise, East Profile" ;
		trise_E:units = "degC" ;
		trise_E:valid_min = 1.f ;
		trise_E:valid_max = 4.5f ;
		trise_E:valid_delta = 3.5f ;
		trise_E:resolution = 0.01f ;
		trise_E:missing_value = -9999.f ;
		trise_E:accuracy = "0.04 degC" ;
	int qc_trise_E(time, depth) ;
		qc_trise_E:long_name = "Quality check results on field: Sensor Temperature Rise, East Profile" ;
		qc_trise_E:units = "unitless" ;
	float soilwatpot_E(time, depth) ;
		soilwatpot_E:long_name = "Soil Water Potential, East Profile" ;
		soilwatpot_E:units = "kPa" ;
		soilwatpot_E:valid_min = -7000.f ;
		soilwatpot_E:valid_max = 0.f ;
		soilwatpot_E:valid_delta = 7000.f ;
		soilwatpot_E:missing_value = -9999.f ;
	int qc_soilwatpot_E(time, depth) ;
		qc_soilwatpot_E:long_name = "Quality check results on field: Soil Water Potential, East Profile" ;
		qc_soilwatpot_E:units = "unitless" ;
	float watcont_E(time, depth) ;
		watcont_E:long_name = "Volumetric Water Content, East Profile" ;
		watcont_E:units = "m3/m3" ;
		watcont_E:valid_min = 0.f ;
		watcont_E:valid_max = 0.55f ;
		watcont_E:valid_delta = 0.55f ;
		watcont_E:missing_value = -9999.f ;
	int qc_watcont_E(time, depth) ;
		qc_watcont_E:long_name = "Quality check results on field: Volumetric Water Content, East Profile" ;
		qc_watcont_E:units = "unitless" ;
	int serial_numbers_W(depth) ;
		serial_numbers_W:long_name = "West profile sensor serial numbers" ;
		serial_numbers_W:units = "unitless" ;
		serial_numbers_W:missing_value = -9999 ;
	int serial_numbers_E(depth) ;
		serial_numbers_E:long_name = "East profile sensor serial numbers" ;
		serial_numbers_E:units = "unitless" ;
		serial_numbers_E:missing_value = -9999 ;
	float lat ;
		lat:long_name = "north latitude" ;
		lat:units = "degrees" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
	float lon ;
		lon:long_name = "east longitude" ;
		lon:units = "degrees" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
	float alt ;
		alt:long_name = "altitude" ;
		alt:units = "meters above Mean Sea Level" ;
	double time(time) ;
		time:units = "seconds since 1970/01/01 00:00:00.00" ;
		time:long_name = "UNIX time" ;

// global attributes:
		:qc_method = "Standard Mentor QC" ;
		:Mentor_QC_Field_Information = "For each qc_<field> interpret the values as follows:\n",
    "\n",
    "Basic mentor QC checks:\n",
    "=======================\n",
    "A value of  0 means that no mentor QC (missing/min/max/delta) checks failed\n",
    "A value of  1 means that the sample contained a \'missing data\' value\n",
    "A value of  2 means that the sample failed the \'minimum\' check\n",
    "A value of  4 means that the sample failed the \'maximum\' check\n",
    "A value of  8 means that the sample failed the \'delta\' check\n",
    "\n",
    "  Note that the delta computation for multi-dimensioned data \n",
    "  compares the absolute value between points in the same spatial \n",
    "  location, at the next point in time. \n",
    "\n",
    "Possible Combinations of mentor QC check results:\n",
    "=================================================\n",
    "\n",
    "A value of  3 means that the sample failed the \'missing and minimum\' checks\n",
    "A value of  5 means that the sample failed the \'missing and maximum\' checks\n",
    "A value of  7 means that the sample failed the \'missing, minimum and maximum\' checks\n",
    "A value of  9 means that the sample failed the \'missing and delta\' checks\n",
    "A value of 10 means that the sample failed the \'minimum and delta\' checks\n",
    "A value of 11 means that the sample failed the \'missing, minimum and delta\' checks\n",
    "A value of 12 means that the sample failed the \'maximum and delta\' checks\n",
    "A value of 14 means that the sample failed the \'minimum, maximum and delta\' checks\n",
    "A value of 15 means that the sample failed the \'missing, minimum, maximum and delta\' checks\n",
    "\n",
    "If the associated non-QC field does not contain any mentor-specified minimum,\n",
    "maximum or delta information, we do not generate a qc_field.\n",
    "" ;
		:mqc_software = "$Id$" ;
		:proc_level = "b1" ;
		:ingest_software = " swats_ingest.c,v 7.2 2001/08/08 04:59:19 ermold process-ingest-swats_ingest-7.4-0 $" ;
		:input_source = "a1 file generated from: swats13:/data/collection/sgp/sgpswatsE13.00/1051747620.icm" ;
		:site_id = "sgp" ;
		:facility_id = "E13 : Lamont_CF1" ;
		:sample_int = "1 hour" ;
		:averaging_int = "not averaged" ;
		:serial_number = "See serial_number data for East and West profiles" ;
		:comment = " " ;
		:resolution_description = "The resolution field attributes refer to the number of significant\n",
    "digits relative to the decimal point that should be used in\n",
    "calculations.  Using fewer digits might result in greater uncertainty;\n",
    "using a larger number of digits should have no effect and thus is\n",
    "unnecessary.  However, analyses based on differences in values with\n",
    "a larger number of significant digits than indicated could lead to\n",
    "erroneous results or misleading scientific conclusions.\n",
    "\n",
    "resolution for lat= 0.001\n",
    "resolution for lon = 0.001\n",
    "resolution for alt = 1" ;
		:profile_distance = "1.0 meter between East and West sensor profiles." ;
		:ref_therm_location = "The reference thermistor is located inside the electronics enclosure which is\n",
    "mounted on a concrete pad sitting on the soil surface. That makes it 1.2m south\n",
    "of the two sensor profiles and 15 cm above the soil surface." ;
		:unit_comment = "kPa is kilopascals, m3/m3 is cubic meters of water per cubic meter of soil." ;
		:soil_characterization = "E13 (Central Facility) This site is located on a broad hilltop, with the\n",
    "topmost sandstone layer about 88 cm below the surface. SWATS sensors are\n",
    "installed at depths of 5, 15, 25, 35, 60, and 85 cm in both profiles.\n",
    "Note: the original installation in late January, 1996 only included the top\n",
    "five levels. The lowest depth (85 cm) was added on 28 February 1997.\n",
    "\n",
    "West 5cm    silt-loam\n",
    "West 15cm   silt-loam\n",
    "West 25cm   clay\n",
    "West 35cm   clay-loam\n",
    "West 60cm   clay-loam\n",
    "West 85cm   clay-loam\n",
    "West 125cm  n/a\n",
    "West 175cm  n/a\n",
    "East 5cm    silt-loam\n",
    "East 15cm   silt-loam\n",
    "East 25cm   clay\n",
    "East 35cm   clay-loam\n",
    "East 60cm   clay-loam\n",
    "East 85cm   clay-loam\n",
    "East 125cm  n/a\n",
    "East 175cm  n/a" ;
		:calib_description = "Calibration/Calculation Technique for determining Soil Water Potential and\n",
    "Volumetric Water Content from the measured SWATS temperature rise values.\n",
    "\n",
    "  Adjustment of individual sensor responses to the \"reference\" sensor response\n",
    "  to remove sensor-to-sensor variability. Coefficients m and b are unique for\n",
    "  each individual sensor.\n",
    "\n",
    "      dTref = m * dTsensor + b\n",
    "\n",
    "    where:\n",
    "\n",
    "      dTref    = \"reference\" sensor response (degC)\n",
    "      dTsensor = individual sensor response  (degC)\n",
    "      m        = slope\n",
    "      b        = intercept\n",
    "\n",
    "    Note: The dTsensor value is input from the \'trise\' fields as reported by\n",
    "    the instrument. However, the dTref value calculated here is NOT the value\n",
    "    stored in the \'tref\' field. This dTref value is only used in the\n",
    "    following calculation.\n",
    "\n",
    "  Second generation calibration used to calculate the soil water potential.\n",
    "\n",
    "      psi = -c * exp(a * dTref)\n",
    "\n",
    "    where:\n",
    "\n",
    "      psi = soil water potential (kPa)\n",
    "      a   = 1.788\n",
    "      c   = 0.717\n",
    "\n",
    "    Note: The value stored in the \'soilwatpot\' field is psi.\n",
    "\n",
    "  Second generation calibration for estimating the water content as a function\n",
    "  of potential. Coefficients tr, ts, alpha, and n are unique for each different\n",
    "  soil layer at each site.\n",
    "\n",
    "      theta = tr + (ts - tr)/(1 + (alpha * (-psi/100))^n)^(1 - 1/n)\n",
    "\n",
    "    where:\n",
    "\n",
    "      theta = volumetric soil water content (m3/m3)\n",
    "      tr    = residual water content (m3/m3)\n",
    "      ts    = saturated water content (m3/m3)\n",
    "      alpha = empirical constant\n",
    "      n     = empirical constant\n",
    "      psi   = potential (kPa)\n",
    "\n",
    "    Note: The value stored in the \'watcont\' field is theta." ;
		:calib_coeficients = "loc\t   m\t   b\t   tr\t   ts\t alpha\t   n\n",
    "w5\t 1.036\t-0.320\t 0.246\t 0.434\t 29.910\t 1.631\n",
    "w15\t 0.990\t-0.244\t 0.246\t 0.434\t 29.910\t 1.631\n",
    "w25\t 1.059\t-0.378\t 0.265\t 0.483\t 66.002\t 1.524\n",
    "w35\t 1.003\t-0.145\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "w60\t 0.950\t-0.159\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "w85\t 1.097\t-0.639\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "w125\t-9999\t-9999\t-9999\t-9999\t-9999\t-9999\n",
    "w175\t-9999\t-9999\t-9999\t-9999\t-9999\t-9999\n",
    "e5\t 1.258\t-0.671\t 0.246\t 0.434\t 29.910\t 1.631\n",
    "e15\t 1.084\t-0.279\t 0.246\t 0.434\t 29.910\t 1.631\n",
    "e25\t 1.044\t-0.354\t 0.265\t 0.483\t 66.002\t 1.524\n",
    "e35\t 1.061\t-0.201\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "e60\t 1.081\t-0.328\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "e85\t 1.071\t 0.073\t 0.297\t 0.479\t 92.101\t 1.284\n",
    "e125\t-9999\t-9999\t-9999\t-9999\t-9999\t-9999\n",
    "e175\t-9999\t-9999\t-9999\t-9999\t-9999\t-9999\n",
    "" ;
		:zeb_platform = "sgpswatsE13.b1" ;
		:history = "Tue Dec  6 06:36:59 2005: ncrcat added variable time=base_time+time_offset\n",
    "Tue Dec  6 06:36:59 2005: ncrcat sgpswatsE13.b1.20030501.000700.cdf sgpswatsE13.b1.20030502.000700.cdf sgpswatsE13.b1.20030503.000700.cdf sgpswatsE13.b1.20030504.000700.cdf sgpswatsE13.b1.20030505.000700.cdf sgpswatsE13.b1.20030506.000700.cdf sgpswatsE13.b1.20030507.000700.cdf sgpswatsE13.b1.20030508.000700.cdf sgpswatsE13.b1.20030509.000700.cdf sgpswatsE13.b1.20030510.000700.cdf sgpswatsE13.b1.20030511.000700.cdf sgpswatsE13.b1.20030512.000700.cdf sgpswatsE13.b1.20030513.000700.cdf sgpswatsE13.b1.20030514.000700.cdf sgpswatsE13.b1.20030515.000700.cdf sgpswatsE13.b1.20030516.000700.cdf sgpswatsE13.b1.20030517.000700.cdf sgpswatsE13.b1.20030518.000700.cdf sgpswatsE13.b1.20030519.000700.cdf sgpswatsE13.b1.20030520.000700.cdf sgpswatsE13.b1.20030521.000700.cdf sgpswatsE13.b1.20030522.000700.cdf sgpswatsE13.b1.20030523.000700.cdf sgpswatsE13.b1.20030524.000700.cdf sgpswatsE13.b1.20030525.000700.cdf sgpswatsE13.b1.20030526.000700.cdf sgpswatsE13.b1.20030527.000700.cdf sgpswatsE13.b1.20030528.000700.cdf sgpswatsE13.b1.20030529.000700.cdf sgpswatsE13.b1.20030530.000700.cdf sgpswatsE13.b1.20030531.000700.cdf sgpswatsE13.b1.20030601.000700.cdf sgpswatsE13.b1.20030602.000700.cdf sgpswatsE13.b1.20030603.000700.cdf sgpswatsE13.b1.20030604.000700.cdf sgpswatsE13.b1.20030605.000700.cdf sgpswatsE13.b1.20030606.000700.cdf sgpswatsE13.b1.20030607.000700.cdf sgpswatsE13.b1.20030608.000700.cdf sgpswatsE13.b1.20030609.000700.cdf sgpswatsE13.b1.20030610.000700.cdf sgpswatsE13.b1.20030611.000700.cdf sgpswatsE13.b1.20030612.000700.cdf sgpswatsE13.b1.20030613.000700.cdf sgpswatsE13.b1.20030614.000700.cdf sgpswatsE13.b1.20030615.000700.cdf sgpswatsE13.b1.20030616.000700.cdf sgpswatsE13.b1.20030617.000700.cdf sgpswatsE13.b1.20030618.000700.cdf sgpswatsE13.b1.20030619.000700.cdf sgpswatsE13.b1.20030620.000700.cdf sgpswatsE13.b1.20030621.000700.cdf sgpswatsE13.b1.20030622.000700.cdf sgpswatsE13.b1.20030623.000700.cdf sgpswatsE13.b1.20030624.000700.cdf sgpswatsE13.b1.20030625.000700.cdf sgpswatsE13.b1.20030626.000700.cdf sgpswatsE13.b1.20030627.000700.cdf sgpswatsE13.b1.20030628.000700.cdf sgpswatsE13.b1.20030629.000700.cdf sgpswatsE13.b1.20030630.000700.cdf sgpswatsE13.b1.20030701.000700.cdf sgpswatsE13.b1.20030702.000700.cdf sgpswatsE13.b1.20030703.000700.cdf sgpswatsE13.b1.20030704.000700.cdf sgpswatsE13.b1.20030705.000700.cdf sgpswatsE13.b1.20030706.000700.cdf sgpswatsE13.b1.20030707.000700.cdf sgpswatsE13.b1.20030708.000700.cdf sgpswatsE13.b1.20030709.000700.cdf sgpswatsE13.b1.20030710.000700.cdf sgpswatsE13.b1.20030711.000700.cdf sgpswatsE13.b1.20030712.000700.cdf sgpswatsE13.b1.20030713.000700.cdf sgpswatsE13.b1.20030714.000700.cdf sgpswatsE13.b1.20030715.000700.cdf sgpswatsE13.b1.BAMEX.nc\n",
    "created by user dsmgr on machine left at 1-May-2003,4:39:59, using $State$" ;
}
