netcdf filter_input_diurnal {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 10 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double concentration(time, member, location) ;
		concentration:long_name = "tracer concentration" ;
		concentration:units = "mass" ;

	double mean_source(time, member, location) ;
		mean_source:long_name = "mean source" ;
		mean_source:units = "mass/timestep" ;

	double source(time, member, location) ;
		source:long_name = "source" ;
		source:units = "mass/timestep" ;

	double source_phase(time, member, location) ;
		source_phase:long_name = "source phase" ;
		source_phase:units = "radians" ;

	double wind(time, member, location) ;
		wind:long_name = "wind" ;
		wind:units = "gridpoints/timestep" ;

	double concentration_priorinf_mean(time, location) ;
		concentration_priorinf_mean:long_name = "prior inflation value for concentration" ;

	double mean_source_priorinf_mean(time, location) ;
		mean_source_priorinf_mean:long_name = "prior inflation value for mean source" ;

	double source_phase_priorinf_mean(time, location) ;
		source_phase_priorinf_mean:long_name = "prior inflation value for source phase" ;

	double source_priorinf_mean(time, location) ;
		source_priorinf_mean:long_name = "prior inflation value for source" ;

	double wind_priorinf_mean(time, location) ;
		wind_priorinf_mean:long_name = "prior inflation value for wind" ;

	double concentration_priorinf_sd(time, location) ;
		concentration_priorinf_sd:long_name = "prior inflation standard deviation for concentration" ;

	double mean_source_priorinf_sd(time, location) ;
		mean_source_priorinf_sd:long_name = "prior inflation standard deviation for mean source" ;

	double source_phase_priorinf_sd(time, location) ;
		source_phase_priorinf_sd:long_name = "prior inflation standard deviation for source phase" ;

	double source_priorinf_sd(time, location) ;
		source_priorinf_sd:long_name = "prior inflation standard deviation for source" ;

	double wind_priorinf_sd(time, location) ;
		wind_priorinf_sd:long_name = "prior inflation standard deviation for wind" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;
		location:axis = "X" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
                time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		time:units = "days since 0000-01-01 00:00:00" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "no calendar" ;
		advance_to_time:units = "days since 0000-00-00 00:00:00" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
		:description = "Initial conditions for diurnal cycle in source model" ;
		:model = "simple_advection" ;
		:destruction_rate = 5.555556e-05 ;
		:history = "same values as in filter_ics r3005 (circa July 2007)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 concentration =
  4546.42683149932, 3972.19995226801, 3309.51540303994, 2932.63582201194, 
    2640.05427740856, 2320.14594988783, 2153.3549966327, 1983.52093393512, 
    1805.46712562517, 1706.75613097564,
  4446.68988685287, 3988.86934205587, 3363.31067894392, 2916.42788197581, 
    2633.09211507771, 2333.96196008349, 2189.6402223906, 1972.16790865866, 
    1790.60086236786, 1731.41686016394,
  4535.89292258479, 3984.503396665, 3321.84407196193, 2977.70289481441, 
    2611.11605051325, 2329.70033045295, 2157.170586184, 1949.67631309324, 
    1770.51228552432, 1714.87530283119,
  4504.03375608158, 3998.59538173256, 3309.82641470028, 2920.02355218793, 
    2642.47127209109, 2402.5082433985, 2178.9407357851, 1951.75777822458, 
    1819.48270953915, 1706.36028613896,
  4586.12416775589, 3899.38569391252, 3332.60587652856, 2994.260839346, 
    2725.38229780055, 2367.82779215721, 2155.55190945801, 1983.79886913181, 
    1790.87107835847, 1715.5357882721,
  4439.23968977203, 3883.6739664951, 3332.34119469016, 3003.45124224231, 
    2630.41416450965, 2337.20544795703, 2123.82142947861, 1934.02058265566, 
    1794.07501200067, 1693.62133918848,
  4498.29703402743, 3963.21253661461, 3375.06894142843, 2934.77944939377, 
    2636.04074541068, 2351.31121145143, 2142.54734506974, 1996.77060167731, 
    1782.92207870557, 1700.47281609793,
  4572.06219445592, 3940.6887079051, 3309.90896664612, 2924.34893811791, 
    2584.05097258422, 2330.19152542715, 2163.17412241129, 1970.01469100591, 
    1823.98468479309, 1708.746210376,
  4539.76663544292, 3911.47381186535, 3383.41218152329, 2939.99101093864, 
    2641.83617949051, 2316.50303767901, 2196.98677688392, 1986.19747031961, 
    1798.28153320056, 1694.0901386826,
  4412.7549532356, 3920.33697993763, 3392.63174316731, 2937.99078362835, 
    2597.07687072564, 2328.73397006858, 2128.3278460597, 1979.55122075781, 
    1814.06994881892, 1685.10897695131,
  4522.63809997819, 3926.61287175122, 3299.18851126821, 2938.96416100808, 
    2606.30313595692, 2352.2231691533, 2182.50722229597, 1990.2767495291, 
    1799.95542132202, 1679.65331941286,
  4512.50407927512, 3984.20496896034, 3343.58221103605, 2984.35728311989, 
    2627.56878339274, 2321.22826695565, 2121.52991133634, 2004.25627629835, 
    1778.40384211529, 1694.8144062224,
  4498.75654086148, 3944.64082086536, 3347.02036450797, 2961.59409883925, 
    2636.8772174749, 2349.99005340106, 2149.79440545499, 1973.25728517395, 
    1784.48915402531, 1722.33794815004,
  4538.65844440224, 3909.42317173294, 3345.48505930937, 2956.19325823296, 
    2593.06102618223, 2391.58019976035, 2152.5932472773, 1943.99186363959, 
    1813.73288596464, 1681.56776683853,
  4510.75963491909, 3988.53207159507, 3332.02980017479, 3016.5031000871, 
    2586.31907760358, 2367.02864856385, 2148.92716729652, 1949.31663826148, 
    1844.60617873271, 1702.92208225261,
  4535.37969970894, 3955.86664267907, 3314.29457449726, 2992.98672272417, 
    2616.92035362922, 2336.29984699437, 2136.91535306808, 1970.77156790322, 
    1797.45649315011, 1708.31067694274,
  4543.31850155928, 3955.93520088496, 3382.51277465646, 2951.88359902794, 
    2647.02578863856, 2334.90879776801, 2139.01997754598, 2013.25450598392, 
    1822.80736182924, 1715.27128379932,
  4445.38885377101, 3954.45465786233, 3294.2828273209, 2908.02997469917, 
    2623.52815054416, 2341.40514974138, 2143.51425605202, 1972.61356945519, 
    1788.87535473667, 1724.3722209794,
  4461.10530365487, 3969.96073952646, 3307.172524332, 2945.48178587927, 
    2652.04930392459, 2344.5719840301, 2165.43810565341, 1958.42033927085, 
    1789.67775526203, 1702.87783726253,
  4512.50006299547, 3950.14257155067, 3405.6341785851, 2926.81186390697, 
    2665.39803473874, 2367.58739539473, 2127.42015600072, 1954.52815459684, 
    1812.38981001257, 1713.07411656148,
  4550.22124697173, 3923.79799382201, 3346.59483758998, 2943.42862984204, 
    2644.88713091593, 2350.74943506181, 2146.99161609715, 1965.27563701833, 
    1758.00722816139, 1692.7043276265,
  4544.02875940155, 3918.88678706754, 3325.86558361138, 2976.4050440364, 
    2596.16680247678, 2372.74866809169, 2160.38890281003, 1968.50807952941, 
    1794.70299809031, 1703.97482072079,
  4423.41291928019, 3981.07617840227, 3328.03667556029, 2973.86678794174, 
    2651.29748491192, 2327.67187478324, 2142.82070120458, 1985.41879817609, 
    1794.61859413369, 1693.14545045278,
  4463.33134744403, 3929.89221956003, 3392.27390046462, 2870.36971389573, 
    2631.00488243709, 2365.63642537319, 2122.57677512035, 1954.68136647684, 
    1810.20255387364, 1721.97631271275,
  4459.16831018046, 3948.71886095649, 3319.87785087544, 2954.81594685219, 
    2632.95590541664, 2380.04221785707, 2143.88222827607, 1959.60489350088, 
    1795.96963944882, 1713.22737485985,
  4475.76361452358, 3981.10130866083, 3327.60851616973, 2940.16401103405, 
    2640.31014113039, 2343.58484143954, 2146.18690620269, 1971.05885963259, 
    1823.62795308743, 1751.08515912771,
  4530.20087794184, 3912.3867272386, 3348.71437443116, 2938.99015135181, 
    2605.38524274372, 2346.95166920535, 2131.16623568789, 1976.87636462226, 
    1830.22266744424, 1732.54974044262,
  4486.20557502904, 3929.96738501919, 3301.08793876475, 3007.97507073406, 
    2641.58560300604, 2334.6720291844, 2117.594783958, 1985.89508675283, 
    1801.61460742186, 1726.42306570752,
  4496.53114704927, 3934.96782668387, 3311.18094397773, 2955.57201465309, 
    2667.3429559297, 2325.26036205874, 2147.18684881906, 1941.87123318851, 
    1799.1000086573, 1692.85357538424,
  4523.77767851825, 3934.48091080421, 3347.73208692271, 2940.91028260852, 
    2650.50782972158, 2361.39524706686, 2144.73406421029, 1996.9134941359, 
    1824.84018616637, 1700.60634356537,
  4422.70040479527, 3922.11443441216, 3310.69725880157, 2976.31828601456, 
    2618.65743538744, 2341.00385130056, 2143.9385271743, 1986.32202930541, 
    1804.59584863627, 1717.62753630449,
  4448.48275618612, 3995.42951155523, 3320.16139019568, 2933.88282004724, 
    2673.45244763063, 2376.85197190545, 2146.79350346374, 1965.53039657929, 
    1837.5507653673, 1731.72469141608,
  4512.45402747137, 3844.2316538198, 3317.20365584023, 2907.09530559057, 
    2639.76412003192, 2316.526660854, 2182.52532198249, 1968.69132952155, 
    1802.04633323131, 1726.19755090173,
  4450.91573047888, 3940.47725183693, 3296.78172999221, 2956.75417658104, 
    2607.55520014338, 2369.51094489494, 2153.45724096404, 1957.80252419702, 
    1797.91965618568, 1714.34935003665,
  4489.53349529024, 3947.75239903568, 3340.06290826133, 2925.09240162733, 
    2626.2759977003, 2392.91102527947, 2143.67942381187, 1966.3650760846, 
    1800.91437535303, 1704.76173008177,
  4404.27684784347, 3951.64877969714, 3337.54192292352, 2909.51910743185, 
    2595.28387565632, 2340.75536361901, 2135.37063404157, 1970.06279275929, 
    1801.18684688618, 1710.10518608231,
  4465.80055270081, 3969.64230755926, 3360.47830539323, 2992.73838848272, 
    2621.89402694769, 2368.49593501247, 2131.92019086186, 1965.89706387673, 
    1810.82086962663, 1724.76294955805,
  4452.80631506399, 3946.61479965141, 3314.46162946768, 2926.38490257744, 
    2642.88681420208, 2374.75924181268, 2140.75546088494, 1980.38929500644, 
    1812.84915179889, 1728.0409349225,
  4542.52092513046, 3937.00180535762, 3376.06335595571, 2932.72429613976, 
    2613.67602730318, 2380.02305712904, 2119.27618342241, 1917.7027168613, 
    1810.26825465819, 1714.0183222836,
  4459.17287817487, 3953.61703426473, 3393.30648760084, 2969.98517274028, 
    2635.49599171277, 2322.49710884252, 2169.76987724974, 1958.63229785199, 
    1798.74230305936, 1709.34962904978,
  4495.58702893491, 3980.64101668237, 3403.10168824038, 2919.56020217178, 
    2650.91924920269, 2351.58034761275, 2153.7553532506, 1977.11787585759, 
    1776.29558654235, 1705.50038793249,
  4428.38910696222, 3963.23165285124, 3311.36813746375, 2942.47360482965, 
    2618.25262446308, 2377.09225762998, 2176.40223872724, 1977.52839859546, 
    1800.85180328687, 1716.29619352612,
  4476.87280589795, 3948.12713711015, 3329.35494685443, 2941.50395158183, 
    2685.43684332057, 2366.96528558965, 2139.54675606331, 1945.5705322332, 
    1797.18922257337, 1694.11650032024,
  4490.81369437315, 3931.42253654618, 3343.42343674938, 2946.48569515356, 
    2669.21702253885, 2321.75938485885, 2159.54075341613, 1948.77386314907, 
    1821.08001253696, 1712.15943446224,
  4511.90117009531, 3934.00862492237, 3343.7549448576, 2957.11132741493, 
    2613.72799064092, 2364.56015508979, 2152.14374625567, 1965.06364443176, 
    1799.62722841858, 1723.59360639749,
  4512.9031811218, 3950.28099740619, 3366.3716480719, 2932.81146780291, 
    2634.53270553383, 2321.96161287962, 2160.50420384221, 1975.16918542003, 
    1861.24526803672, 1716.24695706553,
  4558.6910925682, 3936.11452751085, 3272.20882792954, 2977.64437530228, 
    2591.65767389978, 2296.18825277277, 2131.96254134888, 1969.45273987036, 
    1765.88453322662, 1704.03738386457,
  4498.61596829917, 3941.90207792416, 3329.64785930627, 2928.20254730364, 
    2659.12064501796, 2361.60009766852, 2137.81700293946, 1952.12234691425, 
    1787.96152491202, 1693.41355578679,
  4479.50180473856, 3922.90756869055, 3312.04027861334, 2967.68095396939, 
    2610.60929637054, 2377.06715474329, 2183.91425326717, 1975.11925433002, 
    1810.34124682575, 1718.90221368453,
  4457.75380732031, 3991.97655783437, 3301.44621264942, 2957.62967684282, 
    2621.15935337849, 2320.73682615758, 2127.52173235781, 1980.95536935887, 
    1812.19387615944, 1725.4699160726,
  4511.8089160679, 3917.08410506803, 3305.86243884904, 2975.52113243827, 
    2663.02698200195, 2346.32700697778, 2133.6360878561, 1951.93887223238, 
    1812.75583142417, 1746.3957701225,
  4500.49018299373, 3918.38552791372, 3325.76911958198, 2938.87171474829, 
    2565.14276279008, 2373.13190598408, 2152.40998587666, 1969.51996711232, 
    1796.79204349947, 1708.86298736827,
  4519.24911609974, 3934.47032120745, 3333.28145144799, 2938.72605453766, 
    2586.61653629234, 2413.08281359491, 2143.32051824248, 2022.01619423319, 
    1793.13478983626, 1736.24113396401,
  4530.66499225645, 3928.90523885143, 3294.57501693009, 2949.50807690803, 
    2624.47216949877, 2345.35505775898, 2089.64841475974, 1987.75075215866, 
    1825.97396154421, 1712.01911233598,
  4451.59938008639, 3966.0057746334, 3365.20605309802, 2942.7821335533, 
    2621.29450390212, 2351.5805023835, 2179.68560845463, 1956.57673035976, 
    1794.0751798349, 1727.79896511549,
  4554.20474187022, 3954.9662788884, 3358.12806848645, 2961.51697767998, 
    2615.32130836914, 2330.27465804995, 2182.79324048446, 1979.30045964241, 
    1802.2926162062, 1705.83984822771,
  4489.85992037769, 3928.70561813242, 3347.68074589245, 2934.5885511175, 
    2621.97824154627, 2334.38791329674, 2112.34604111985, 1995.55455771731, 
    1787.0474324849, 1705.6410255713,
  4487.09012489022, 3971.49632930666, 3297.81351962914, 2984.42200951886, 
    2619.28706945478, 2372.42349288841, 2163.9386592018, 1948.75180630289, 
    1796.09889875553, 1714.6864488463,
  4465.49289388225, 4001.91670531823, 3329.68475703834, 2910.81970987924, 
    2610.68793449922, 2344.96020494913, 2151.36067655503, 1967.13636361595, 
    1810.02377285551, 1716.41890653485,
  4433.26919926666, 3949.21589912298, 3318.26545151891, 2938.35592794045, 
    2637.90340243797, 2346.4041475625, 2157.25487657919, 1960.15430916486, 
    1796.74716332572, 1705.11616071626,
  4486.26484591613, 3923.2189462125, 3410.51306530546, 2920.74435385744, 
    2660.70664986067, 2336.34011779718, 2150.91669416099, 1957.51874796904, 
    1802.31268280302, 1712.49512004532,
  4499.20321653197, 3923.38055562591, 3384.80524450793, 2991.78762652344, 
    2617.99312781837, 2354.99994434918, 2133.27979041304, 1948.02834356999, 
    1817.60317189196, 1705.72626150919,
  4581.45146499614, 3920.11181902053, 3346.89929602008, 2977.30967651251, 
    2601.08877527274, 2360.50519738454, 2157.60137717075, 1995.48142502575, 
    1794.11682701832, 1689.10517442201,
  4506.2375304021, 3919.162964825, 3339.6006190538, 2890.31387282688, 
    2654.48247321565, 2378.1201415219, 2155.38740595177, 1975.6245722382, 
    1797.66070127017, 1692.82503029414,
  4445.45542915109, 3980.43525395572, 3342.0575985534, 2938.28934429396, 
    2628.29445224313, 2322.6982199671, 2132.00941225448, 1930.81154726013, 
    1780.21383515986, 1716.9695136981,
  4459.3881812794, 3899.99068344037, 3319.33009331264, 2962.14693519106, 
    2663.27303699728, 2306.39837641447, 2144.80817163425, 2003.44586616826, 
    1796.68055729016, 1717.4967836512,
  4591.36035458122, 3934.12428468785, 3317.59391411651, 2937.51007705099, 
    2651.41880140734, 2355.57790400643, 2165.11503053252, 1945.97173114149, 
    1800.87860414671, 1699.22152594411,
  4479.5588598518, 3957.6199255654, 3345.29985549307, 2975.51286254328, 
    2636.6684172735, 2331.19250227739, 2166.16196612834, 1951.16352200635, 
    1793.84526316648, 1714.30103230276,
  4460.48515608559, 3940.88193566056, 3311.46557927438, 2995.50138599886, 
    2625.07806901497, 2352.92363066057, 2145.01620918455, 1953.34739264613, 
    1812.58837681625, 1725.47463468238,
  4369.14116889016, 3989.68714308314, 3334.62249421548, 3036.65947248928, 
    2632.77529740527, 2362.96125620693, 2214.3630277445, 1983.41327283837, 
    1809.46055547826, 1729.74938665808,
  4422.25645548906, 3971.95933780118, 3355.21436514089, 2941.67877135216, 
    2634.52680141934, 2338.50495673667, 2153.86045777987, 1988.24029910136, 
    1802.29696078617, 1707.62953546177,
  4468.99493475593, 3910.33714174466, 3338.52362498405, 2903.16269360897, 
    2695.86410467179, 2363.0635365889, 2133.65247565732, 1945.34515001226, 
    1788.96407042978, 1709.49622102573,
  4534.90574720455, 3970.25003552501, 3312.16104964452, 2953.86958097514, 
    2664.99681252151, 2369.37326810839, 2156.304168164, 1989.55259376013, 
    1800.89406659513, 1710.14995194385,
  4433.16585770015, 3997.83982649106, 3256.12977651173, 2970.02861299539, 
    2596.30234747301, 2382.26887584704, 2145.92721427845, 1974.02524649376, 
    1792.71782927099, 1723.98445330203,
  4550.59585378827, 3934.79148013725, 3328.98378748163, 2917.22001745559, 
    2654.23977494549, 2327.05727869178, 2122.93790441409, 1958.14064060409, 
    1812.62266888372, 1713.92272556888,
  4451.7797253039, 3938.60459407083, 3337.86482210721, 2925.06023292906, 
    2661.1275031082, 2372.01380480406, 2134.63538544532, 2022.52573347979, 
    1839.73860356767, 1700.00757780891,
  4573.60192025348, 3954.6784310962, 3317.14268533638, 2926.34687663542, 
    2650.08860799036, 2357.23577717672, 2143.40268745771, 1959.65657310954, 
    1799.22069853874, 1688.58550781623,
  4483.11932280885, 3964.16082183253, 3337.61242722367, 2951.54933943067, 
    2632.91363425624, 2350.78169363328, 2159.7999484092, 1993.83109639755, 
    1825.84080145668, 1712.8370993246,
  4482.80396847085, 3937.03901256269, 3352.08565747793, 3021.37250490131, 
    2624.52845917467, 2387.34801849286, 2132.47294857178, 1995.50333064304, 
    1815.66116667526, 1721.8621266059,
  4505.17745668008, 3910.97736469217, 3319.32539023918, 2950.73795423536, 
    2634.49616107807, 2314.01198771261, 2159.3766919411, 1971.15818123444, 
    1801.67183752271, 1730.67358960651 ;

 mean_source =
  1.00000000000149, 0.100000000000147, 0.100000000000147, 0.100000000000147, 
    0.100000000000147, 0.100000000000147, 0.100000000000147, 
    0.100000000000147, 0.100000000000147, 0.100000000000147,
  1.00000000000161, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016,
  1.00000000000145, 0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144,
  1.00000000000146, 0.100000000000145, 0.100000000000145, 0.100000000000145, 
    0.100000000000145, 0.100000000000145, 0.100000000000145, 
    0.100000000000145, 0.100000000000145, 0.100000000000145,
  1.00000000000156, 0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155,
  1.00000000000161, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016,
  1.0000000000016, 0.100000000000159, 0.100000000000159, 0.100000000000159, 
    0.100000000000159, 0.100000000000159, 0.100000000000159, 
    0.100000000000159, 0.100000000000159, 0.100000000000159,
  1.0000000000014, 0.100000000000139, 0.100000000000139, 0.100000000000139, 
    0.100000000000139, 0.100000000000139, 0.100000000000139, 
    0.100000000000139, 0.100000000000139, 0.100000000000139,
  1.00000000000159, 0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158,
  1.00000000000164, 0.100000000000163, 0.100000000000163, 0.100000000000163, 
    0.100000000000163, 0.100000000000163, 0.100000000000163, 
    0.100000000000163, 0.100000000000163, 0.100000000000163,
  1.00000000000155, 0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154,
  1.00000000000142, 0.100000000000141, 0.100000000000141, 0.100000000000141, 
    0.100000000000141, 0.100000000000141, 0.100000000000141, 
    0.100000000000141, 0.100000000000141, 0.100000000000141,
  1.0000000000015, 0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149,
  1.0000000000017, 0.100000000000169, 0.100000000000169, 0.100000000000169, 
    0.100000000000169, 0.100000000000169, 0.100000000000169, 
    0.100000000000169, 0.100000000000169, 0.100000000000169,
  1.00000000000149, 0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149,
  1.00000000000156, 0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155,
  1.00000000000165, 0.100000000000164, 0.100000000000164, 0.100000000000164, 
    0.100000000000164, 0.100000000000164, 0.100000000000164, 
    0.100000000000164, 0.100000000000164, 0.100000000000164,
  1.00000000000148, 0.100000000000147, 0.100000000000147, 0.100000000000147, 
    0.100000000000147, 0.100000000000147, 0.100000000000147, 
    0.100000000000147, 0.100000000000147, 0.100000000000147,
  1.00000000000161, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016, 0.10000000000016, 0.10000000000016, 
    0.10000000000016, 0.10000000000016,
  1.00000000000167, 0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166,
  1.00000000000154, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000151, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015,
  1.00000000000144, 0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144,
  1.00000000000156, 0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155,
  1.00000000000141, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014,
  1.00000000000145, 0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144,
  1.00000000000151, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015,
  1.00000000000154, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000159, 0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158,
  1.00000000000155, 0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155,
  1.00000000000142, 0.100000000000141, 0.100000000000141, 0.100000000000141, 
    0.100000000000141, 0.100000000000141, 0.100000000000141, 
    0.100000000000141, 0.100000000000141, 0.100000000000141,
  1.00000000000154, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.0000000000015, 0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149,
  1.00000000000156, 0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155, 
    0.100000000000155, 0.100000000000155, 0.100000000000155,
  1.00000000000157, 0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156,
  1.00000000000155, 0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154,
  1.00000000000152, 0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151,
  1.00000000000141, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014,
  1.00000000000158, 0.100000000000157, 0.100000000000157, 0.100000000000157, 
    0.100000000000157, 0.100000000000157, 0.100000000000157, 
    0.100000000000157, 0.100000000000157, 0.100000000000157,
  1.0000000000015, 0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149,
  1.0000000000016, 0.100000000000159, 0.100000000000159, 0.100000000000159, 
    0.100000000000159, 0.100000000000159, 0.100000000000159, 
    0.100000000000159, 0.100000000000159, 0.100000000000159,
  1.00000000000151, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015,
  1.00000000000144, 0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.00000000000162, 0.100000000000161, 0.100000000000161, 0.100000000000161, 
    0.100000000000161, 0.100000000000161, 0.100000000000161, 
    0.100000000000161, 0.100000000000161, 0.100000000000161,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.00000000000153, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000149, 0.100000000000148, 0.100000000000148, 0.100000000000148, 
    0.100000000000148, 0.100000000000148, 0.100000000000148, 
    0.100000000000148, 0.100000000000148, 0.100000000000148,
  1.00000000000155, 0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.00000000000151, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015,
  1.00000000000167, 0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.00000000000154, 0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154,
  1.00000000000157, 0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156,
  1.00000000000174, 0.100000000000173, 0.100000000000173, 0.100000000000173, 
    0.100000000000173, 0.100000000000173, 0.100000000000173, 
    0.100000000000173, 0.100000000000173, 0.100000000000173,
  1.00000000000154, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000153, 0.100000000000152, 0.100000000000152, 0.100000000000152, 
    0.100000000000152, 0.100000000000152, 0.100000000000152, 
    0.100000000000152, 0.100000000000152, 0.100000000000152,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.0000000000015, 0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149, 
    0.100000000000149, 0.100000000000149, 0.100000000000149,
  1.00000000000155, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000167, 0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166, 
    0.100000000000166, 0.100000000000166, 0.100000000000166,
  1.00000000000155, 0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154, 
    0.100000000000154, 0.100000000000154, 0.100000000000154,
  1.00000000000159, 0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158,
  1.00000000000145, 0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144, 
    0.100000000000144, 0.100000000000144, 0.100000000000144,
  1.00000000000151, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015, 0.10000000000015, 0.10000000000015, 
    0.10000000000015, 0.10000000000015,
  1.00000000000153, 0.100000000000152, 0.100000000000152, 0.100000000000152, 
    0.100000000000152, 0.100000000000152, 0.100000000000152, 
    0.100000000000152, 0.100000000000152, 0.100000000000152,
  1.00000000000147, 0.100000000000145, 0.100000000000145, 0.100000000000145, 
    0.100000000000145, 0.100000000000145, 0.100000000000145, 
    0.100000000000145, 0.100000000000145, 0.100000000000145,
  1.00000000000143, 0.100000000000142, 0.100000000000142, 0.100000000000142, 
    0.100000000000142, 0.100000000000142, 0.100000000000142, 
    0.100000000000142, 0.100000000000142, 0.100000000000142,
  1.00000000000152, 0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151,
  1.00000000000144, 0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143,
  1.00000000000141, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014, 0.10000000000014, 0.10000000000014, 
    0.10000000000014, 0.10000000000014,
  1.00000000000158, 0.100000000000157, 0.100000000000157, 0.100000000000157, 
    0.100000000000157, 0.100000000000157, 0.100000000000157, 
    0.100000000000157, 0.100000000000157, 0.100000000000157,
  1.00000000000169, 0.100000000000168, 0.100000000000168, 0.100000000000168, 
    0.100000000000168, 0.100000000000168, 0.100000000000168, 
    0.100000000000168, 0.100000000000168, 0.100000000000168,
  1.00000000000147, 0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146, 
    0.100000000000146, 0.100000000000146, 0.100000000000146,
  1.00000000000144, 0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143, 
    0.100000000000143, 0.100000000000143, 0.100000000000143,
  1.00000000000154, 0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153, 
    0.100000000000153, 0.100000000000153, 0.100000000000153,
  1.00000000000159, 0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158, 
    0.100000000000158, 0.100000000000158, 0.100000000000158,
  1.00000000000157, 0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156, 
    0.100000000000156, 0.100000000000156, 0.100000000000156,
  1.00000000000152, 0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151, 
    0.100000000000151, 0.100000000000151, 0.100000000000151 ;

 source =
  0.824569222923133, 0.0784316692637661, 0.0728123553430491, 
    0.0860442480535596, 0.0899233875778706, 0.0807436815569396, 
    0.0868307792177679, 0.07571733946983, 0.0855521088728275, 
    0.0880934328792199,
  0.816695618523789, 0.0917850410223096, 0.0706698466840174, 
    0.0875382162438299, 0.0842465778637555, 0.0815055961094878, 
    0.0897114728034078, 0.083823935485998, 0.0860507269868346, 
    0.0901875806199394,
  0.840666802536394, 0.0871971318439315, 0.0727446472054706, 
    0.0940625853373903, 0.0802252087575856, 0.0826256345749374, 
    0.0849075074307129, 0.0825705947857377, 0.07763671495784, 
    0.0950266446720765,
  0.845822666824601, 0.0879586040596868, 0.0764188790540102, 
    0.0924640845091722, 0.0867285162569057, 0.0786260184137855, 
    0.0857231126112958, 0.0790529407584183, 0.0840690230876636, 
    0.0878300759214507,
  0.825745982166528, 0.0893673508453082, 0.0657427363019919, 
    0.0993360786529308, 0.0792637823110335, 0.0889663707948512, 
    0.0878709863195418, 0.0836747684286982, 0.0801714557124375, 
    0.0909608740506254,
  0.80090924191954, 0.0883928328863767, 0.0763459524947668, 
    0.0893941108505044, 0.090178074008068, 0.0836649759060446, 
    0.0843928792056054, 0.0782248145763484, 0.0842977653522912, 
    0.0842094693378455,
  0.828126488857206, 0.0843347922084905, 0.0749536754662669, 
    0.0875533852188562, 0.0898706763296858, 0.0822767649728138, 
    0.083689879380598, 0.0853173456330593, 0.080340280514714, 
    0.0916485753562901,
  0.808321741124625, 0.0889730815130887, 0.0758862320311772, 
    0.0896377101022729, 0.0768929452745882, 0.0838315934627605, 
    0.0839332550581607, 0.0809539028927209, 0.0886014119445543, 
    0.0851966926760962,
  0.848985832714675, 0.0823335164316614, 0.087729589100141, 
    0.0812265111105321, 0.0900815455211044, 0.0795809940646528, 
    0.097131631716846, 0.0771213066610647, 0.0786420805044018, 
    0.090463221813171,
  0.825376823214736, 0.0880098934162369, 0.0781010623041865, 
    0.0880769693309879, 0.0723872579443663, 0.0828281433626209, 
    0.089836524177917, 0.0802604706034371, 0.0880377937702971, 
    0.0827359544415985,
  0.852899857226161, 0.0822638255197437, 0.0764104513815365, 
    0.0945834975791768, 0.0765099198181105, 0.0908929359827314, 
    0.08606464915903, 0.0814149632600218, 0.0782418944355277, 
    0.0880826000200291,
  0.811334379821341, 0.088401818629605, 0.0745250972185029, 
    0.0914639700535213, 0.0759185885900142, 0.0879727308271168, 
    0.0853458192887898, 0.0783769903052301, 0.083660513609383, 
    0.0884207660550121,
  0.841832954953528, 0.0860847483783202, 0.0774423337148951, 
    0.0977767053595035, 0.0710746573893921, 0.0870942657632219, 
    0.0856866507070514, 0.0786600274117655, 0.0783002843862242, 
    0.0953436892444174,
  0.864545641409224, 0.089673199183141, 0.0800891250096354, 
    0.0922151018586243, 0.0745729297239055, 0.0896466134309217, 
    0.0877874807714002, 0.0859929721336801, 0.0811361515371092, 
    0.0853009570704637,
  0.833533308875256, 0.0838255988394539, 0.082574295373474, 
    0.0884138021737063, 0.0797775678913059, 0.0900421021377545, 
    0.0848639411132848, 0.0789999238009393, 0.0837624138168356, 
    0.0850998917284897,
  0.828438856183434, 0.0832994540035071, 0.0783344895177846, 
    0.0986152506760215, 0.0798458358785261, 0.088644289216717, 
    0.0825852686954762, 0.0827792020683466, 0.0870612220182748, 
    0.0894691913537476,
  0.833568674950937, 0.0875940034008963, 0.074318848120459, 
    0.0941308883144478, 0.0830589480619523, 0.0798375250665419, 
    0.0836395417087894, 0.0849016322610666, 0.0853479316888178, 
    0.0845766771519424,
  0.823194793036184, 0.082144751920925, 0.0755997346379119, 
    0.084103753775088, 0.0860230414323392, 0.0782833852504952, 
    0.0854009348294736, 0.0775484356306201, 0.0848866843324875, 
    0.0935785357176507,
  0.803525066355385, 0.0820122490644355, 0.0717971336695247, 
    0.0908099975530424, 0.0821987127341539, 0.0798332232019284, 
    0.0893016056400799, 0.0785947249112255, 0.084402502491762, 
    0.0864381872123786,
  0.820031349282103, 0.0852830058349414, 0.0706337933753045, 
    0.0837940114547668, 0.0774734111203114, 0.0861362514226402, 
    0.0880824897953685, 0.0790654809955941, 0.0833824429105823, 
    0.0921340754474347,
  0.826297471828937, 0.086717991685809, 0.075611387463316, 
    0.0881729914571785, 0.0872374714810876, 0.0856684984239115, 
    0.0815453739741744, 0.0772781789403963, 0.0754030042943033, 
    0.0869371887578209,
  0.841471903687483, 0.0869256741491669, 0.0761770399449724, 
    0.0869375929528625, 0.0791842295186788, 0.0869805637543107, 
    0.0888701801246906, 0.0791628704508645, 0.0876993389069076, 
    0.0885768644405143,
  0.812170872772817, 0.0882694324339774, 0.0663905750957852, 
    0.0933579942004789, 0.0879143502364382, 0.0796324895735926, 
    0.0866510239716202, 0.079380967801986, 0.0833975867324361, 
    0.0911718413015139,
  0.818272669061862, 0.087699754966837, 0.0751176762414525, 
    0.0896476591483001, 0.0843351181304001, 0.0878217255294105, 
    0.0885000207696341, 0.0821852366112777, 0.0798899717019309, 
    0.0882540731101231,
  0.834489080912413, 0.0861510068800036, 0.0759591998067344, 
    0.0916974853867416, 0.0874521443010292, 0.0887295228207036, 
    0.0863611562547902, 0.0795650225880686, 0.0820666292196929, 
    0.0847876361510181,
  0.830032997501602, 0.0844117355073031, 0.0723352911965123, 
    0.0901925840007655, 0.0828199043701857, 0.0862469725902025, 
    0.0884745030158937, 0.07985162072864, 0.0903980088032482, 
    0.091641753895792,
  0.806836514157933, 0.0918599618159149, 0.0777704592661771, 
    0.0914631331568836, 0.0872989834006049, 0.0834425710158154, 
    0.0868470987847333, 0.0829412658931275, 0.0869775763735076, 
    0.090703599457999,
  0.870336469600163, 0.086219104422921, 0.066651090373386, 
    0.0933057800569064, 0.0793274763218805, 0.0779761859231986, 
    0.0830583584671072, 0.0835260320854172, 0.0805022929804514, 
    0.0890340719605608,
  0.798904613483585, 0.0878182529169572, 0.077430818110271, 
    0.0928965233172025, 0.0817233179638871, 0.0807004545748917, 
    0.0897661630183422, 0.0799034023504768, 0.0887613506623904, 
    0.0886146757286244,
  0.831779634528505, 0.0846560776813716, 0.0723103258739772, 
    0.0860456462276937, 0.083144011993218, 0.0869283053637341, 
    0.0853170012946901, 0.0784333460378027, 0.0872441452912708, 
    0.0870532396580271,
  0.821362520846727, 0.0839968812553347, 0.0763224032231107, 
    0.0896901214864734, 0.0820056240004905, 0.0777055914419637, 
    0.093431757495256, 0.0776376723242199, 0.0761596031488464, 
    0.0939056359934546,
  0.800237779915415, 0.0897015792177949, 0.0695490731811666, 
    0.09454775072917, 0.0857245342091019, 0.077041946086549, 
    0.0915018768565468, 0.0765253511141415, 0.0850764807402921, 
    0.0906392431648071,
  0.794862798195074, 0.0851318127789901, 0.072512332106333, 
    0.0923467145602342, 0.0781355861654487, 0.0856744035600605, 
    0.0921292155319738, 0.0743188339815406, 0.0843349683677926, 
    0.0911662813592882,
  0.782828744207989, 0.0896924924110309, 0.0675648738283316, 
    0.0946267674740224, 0.0807777362492993, 0.0868508390700235, 
    0.0859812064460206, 0.0840585802556364, 0.0829089870539731, 
    0.090842025878781,
  0.813951919996239, 0.0885772966566522, 0.0659476644639829, 
    0.0932307907708749, 0.082981523966751, 0.089443307087404, 
    0.0830859470387562, 0.0800365679929171, 0.0816118816780815, 
    0.0919535875971096,
  0.817708101894119, 0.0927441599486021, 0.0682488185772263, 
    0.0960932129980992, 0.0815751847595522, 0.0879003610806895, 
    0.0868402343018331, 0.0815343892615931, 0.0814901532483186, 
    0.0937924711149639,
  0.846329984234003, 0.0827330239347323, 0.0755800595443339, 
    0.088398484721831, 0.0781606633150549, 0.0875556602397347, 
    0.0852191894881418, 0.0797781035681098, 0.085346571111855, 
    0.0921221744329008,
  0.838579166699302, 0.0897357342507066, 0.0761561013595254, 
    0.0909196860178153, 0.0817403392481528, 0.0822509692108274, 
    0.0834634434882253, 0.0817564516735714, 0.087052283608817, 
    0.0918294786260135,
  0.827776386189886, 0.0883567252853157, 0.0662865626091384, 
    0.0915420387277886, 0.0798040948327688, 0.0838731675815869, 
    0.0867530203037342, 0.0770721055000112, 0.0868269534421285, 
    0.090385411742133,
  0.829277337770845, 0.0902329952721942, 0.0693798037761636, 
    0.0875502794518788, 0.0878219950191202, 0.076387131982999, 
    0.0928125352673206, 0.0795609032377843, 0.0809263731142727, 
    0.090636064431794,
  0.84575249157889, 0.0849280923585945, 0.0823430624493593, 
    0.0928494042109447, 0.0869517082475217, 0.0792553416873741, 
    0.0918494882642479, 0.0778120830169321, 0.0826191579953835, 
    0.0931630643131077,
  0.837293972629568, 0.086149566887489, 0.0641542138728477, 
    0.0890675058977376, 0.0823340204173042, 0.0898986319115619, 
    0.0819151183302112, 0.0860438189612508, 0.0892322429757322, 
    0.0895933501023317,
  0.832863597430142, 0.0829208108336731, 0.0830166202962869, 
    0.0871747874564755, 0.0844387199480811, 0.0888461722369248, 
    0.0840244780689674, 0.081458508856818, 0.0843898727093846, 
    0.0877108593581657,
  0.793553750349707, 0.0809578862692568, 0.0824621125802457, 
    0.0941542613752545, 0.0782199051057353, 0.0911343629295461, 
    0.084088106727107, 0.0807291070205356, 0.0914721857009086, 
    0.0840538895222016,
  0.797265910749895, 0.084647512019815, 0.0757069323271163, 
    0.0890713811926921, 0.0815898242654731, 0.0878430711665781, 
    0.0842366885707598, 0.0827025175367064, 0.0848036972658764, 
    0.0889218842160984,
  0.844668833271491, 0.0876802012761761, 0.0804177399353157, 
    0.0903986248184358, 0.0854204343056674, 0.0788938822820796, 
    0.0896235517980078, 0.0780220273639436, 0.0908666812474734, 
    0.0857694412118815,
  0.858119007809378, 0.0914926545993508, 0.0721045432542372, 
    0.0938960492933803, 0.0802992635432757, 0.082523221592548, 
    0.0875174031623939, 0.0834839093363108, 0.0778811795848136, 
    0.0891993209558969,
  0.840895377467152, 0.0774612441034231, 0.0820298616823118, 
    0.0829002384165858, 0.0837221683858367, 0.0838373595869285, 
    0.0885894951565719, 0.0768485039492269, 0.0826497963403641, 
    0.0850005935802425,
  0.781897501354461, 0.0853353734205984, 0.0740542233220466, 
    0.0910298697764406, 0.0831889476447203, 0.0839950734495294, 
    0.0865146114768722, 0.0756178981215846, 0.0820475659413796, 
    0.0888980663663489,
  0.820053024362188, 0.0855880471214074, 0.0720869003704529, 
    0.0917085317294082, 0.0854400773404779, 0.0825913358322986, 
    0.0827859487166747, 0.0806786552811666, 0.0826034616622051, 
    0.0929193780846374,
  0.814870541454436, 0.0914447182064527, 0.0695200475822885, 
    0.0883331326585186, 0.0841739166385681, 0.082857372445697, 
    0.0885051413011368, 0.0853062872182852, 0.0846024861872689, 
    0.0919867721624555,
  0.84788932650228, 0.0851962693089627, 0.0744231688335327, 
    0.0897927425725246, 0.0779243065001275, 0.083317445639292, 
    0.0818465444653485, 0.0790097973863497, 0.0818030009317825, 
    0.0891345655809971,
  0.832873289918919, 0.085086851732315, 0.0724230302373672, 
    0.0938330015761602, 0.0745274248065442, 0.0933184088978593, 
    0.0827625493195679, 0.0830198619491928, 0.080611665017438, 
    0.0920835054699992,
  0.855769247978261, 0.0828397991130558, 0.0653719182618587, 
    0.0912975934163771, 0.0805472960813101, 0.0841676911548288, 
    0.0800445613589202, 0.086447466291461, 0.0803208644010065, 
    0.0891036380639183,
  0.876163782864482, 0.083754990453414, 0.0755270083270152, 
    0.0984525938233558, 0.0791860000181132, 0.0868141098518735, 
    0.0838110906566402, 0.0795515797041376, 0.0801566544432354, 
    0.0866446157078153,
  0.818744314029311, 0.0931311844224582, 0.0703268885095147, 
    0.088122248610481, 0.0851068379225477, 0.0846877824956252, 
    0.0941177931945639, 0.0802207132389739, 0.081665460057162, 
    0.0923201665855992,
  0.801142993196111, 0.0843080449763135, 0.0701223139869373, 
    0.0944907540518007, 0.0745328775539726, 0.0884140527369024, 
    0.0814744010158331, 0.0835371043004935, 0.0759420853197305, 
    0.093071524005167,
  0.824676823450223, 0.084714567799768, 0.0723988274287743, 
    0.0899966132544863, 0.0767500221153561, 0.0862092672990935, 
    0.0936564714323815, 0.0828440514034913, 0.0828865889461632, 
    0.0909235482137578,
  0.80624557477616, 0.0883141362864402, 0.0809172366864952, 
    0.0892659412024326, 0.0838763379349008, 0.0875190247099807, 
    0.0879209997120701, 0.0836786648949949, 0.0872843539885507, 
    0.0859598344809173,
  0.820232017388411, 0.0871886779611386, 0.0762060821408516, 
    0.0899955624965411, 0.0794818527983197, 0.0841422717297862, 
    0.0853473893983749, 0.0823793054897134, 0.0852106806934801, 
    0.0864397373592465,
  0.834604912108566, 0.0865693252976112, 0.0786414224703611, 
    0.0890714726465222, 0.0864591113573971, 0.0861350963698844, 
    0.0854298548505428, 0.0754617826595733, 0.083153670503659, 
    0.0841831827395778,
  0.854536569500517, 0.0864348428439755, 0.0717631325042199, 
    0.0967571424074896, 0.091740490435227, 0.0830957400118934, 
    0.0862460520061533, 0.0779033696248233, 0.0879465918029253, 
    0.084802113413615,
  0.820473598065396, 0.0839060132525636, 0.0653750719119022, 
    0.0923328681971745, 0.0846681848828238, 0.0811193890040111, 
    0.0910302784285897, 0.0785781384466231, 0.0868505809427945, 
    0.0822333725946763,
  0.846184242010634, 0.0873929348864528, 0.0721655717618542, 
    0.0865320084499257, 0.0872407191361668, 0.0893016234997508, 
    0.0838357616981762, 0.083605670675531, 0.0807411677991229, 
    0.0881099380661831,
  0.848004632331681, 0.0832123685195912, 0.0722475747937363, 
    0.0961509785980645, 0.0865376544112876, 0.0829853595087137, 
    0.0858245702341455, 0.0783945251723962, 0.0857582365788027, 
    0.0907476213941789,
  0.819337021783024, 0.0838557557905962, 0.0816647492363733, 
    0.0926793812432426, 0.0829067426928643, 0.0796072837250854, 
    0.0892624722061718, 0.0815952783781531, 0.0853462168639405, 
    0.0869097729225042,
  0.835544647763767, 0.0841012030375932, 0.078048538522798, 
    0.0944619996041883, 0.0877303876931569, 0.0851127685289967, 
    0.0920014122789325, 0.0779997773305374, 0.0829293979312376, 
    0.0901678997502998,
  0.823277931298135, 0.089664340518521, 0.0867517262370124, 
    0.0939327051227788, 0.0789869344697865, 0.0920937310604096, 
    0.0854146946535459, 0.0816859080333289, 0.0835625691566347, 
    0.090392372120669,
  0.820163657116834, 0.0841121842059976, 0.0822772738965122, 
    0.0833655542336643, 0.0944294981084749, 0.0771368506270274, 
    0.0895462761778126, 0.0817765789053546, 0.0860421998381361, 
    0.0913410034563562,
  0.849502643460341, 0.086138297800296, 0.0708944700308293, 
    0.0962451880250238, 0.0823529026651439, 0.0881274434037799, 
    0.0866568602935915, 0.0810484836042088, 0.0839314284246951, 
    0.0919146878063078,
  0.82736668917435, 0.0880978873762274, 0.0629567038915573, 
    0.0869741450835326, 0.0789795699773215, 0.0817202193338855, 
    0.0877822181316683, 0.0839352805258649, 0.0795883769007203, 
    0.0892734909047991,
  0.821193749763778, 0.0845258435456795, 0.0723537787149763, 
    0.0922838232078134, 0.0893791506679929, 0.08385988508442, 
    0.0913335299073617, 0.0766027795298385, 0.0825843520365481, 
    0.0886011163667249,
  0.794902181039964, 0.0842722716733675, 0.07283730228754, 
    0.0852203772906117, 0.0864781825228675, 0.0751495375660241, 
    0.086581814066448, 0.0794398879767707, 0.0857781541226497, 
    0.0881639728161998,
  0.830328972246274, 0.0862799719755862, 0.0639611209237379, 
    0.0961977021674697, 0.0724847083859218, 0.0917151281363832, 
    0.084222913453178, 0.080251251687565, 0.0801042158237093, 
    0.0877923396715901,
  0.813640263725447, 0.0866364434216728, 0.0743786486646491, 
    0.0899202667588293, 0.0876506987556083, 0.0762931200772289, 
    0.0907583412165206, 0.0829093579616112, 0.0833190155960973, 
    0.0901381197114414,
  0.797271471705744, 0.0848408415830504, 0.0806895364867578, 
    0.0911084571776759, 0.0869152622008114, 0.0856933070586302, 
    0.087783402049676, 0.0830022646870148, 0.0848783620753296, 
    0.0874757190123662,
  0.827882396221416, 0.091689756261262, 0.0698821460980115, 
    0.0902461070759427, 0.0851614628083386, 0.0855990089145921, 
    0.08816196190905, 0.0797743718443202, 0.0830849525120327, 
    0.0865862931852523,
  0.815530762115135, 0.0901780402344337, 0.0818636855725555, 
    0.0844562194433103, 0.0819195281510827, 0.0865061865763209, 
    0.0908139570582054, 0.0829893498673085, 0.0811446507935365, 
    0.08585495096857,
  0.804934272785749, 0.088436237820877, 0.084099459220167, 
    0.0990609420045685, 0.0794068739242336, 0.0902831083136275, 
    0.0828894196476489, 0.0832459275759689, 0.0860731933667122, 
    0.0876544052522991,
  0.788121458128012, 0.0850069471882671, 0.0756848604347252, 
    0.0882593725244297, 0.0888809989559672, 0.0769669608418673, 
    0.0945072617261523, 0.0823183406220398, 0.0820446439285289, 
    0.0917374705061113 ;

 source_phase =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wind =
  19.6251329612142, 21.2251473584064, 19.2697866825434, 20.8862066546423, 
    25.0075035774869, 23.5965658207201, 18.6815006904928, 20.7082955002016, 
    24.8681689728539, 18.93938650335,
  26.0266822153012, 22.6108928016386, 21.8281914863617, 23.3001243932279, 
    25.656041029576, 23.6881651714965, 21.538363958747, 22.5567015206733, 
    23.4241184151587, 22.7102143759513,
  20.1786597337347, 24.1074007585505, 18.3459557623814, 19.7207984059654, 
    23.2984677057012, 20.5438855436312, 20.4248471744194, 23.6226220193981, 
    20.1216201086112, 18.8686849292496,
  20.7588801731395, 22.5935308983057, 20.3262036582563, 19.0918120688107, 
    24.3022765426886, 24.493444148302, 24.8364124609087, 23.9508678278979, 
    23.5767799808986, 23.8906128588746,
  22.0900442651818, 18.4641540423292, 19.5406922944695, 20.9773798158111, 
    22.4487781752671, 25.4515756667045, 20.6052366007707, 21.0800434485375, 
    22.0593976797873, 20.4516479627432,
  23.0092896930431, 19.498330530569, 20.001281743043, 22.2944876012735, 
    26.4532226887918, 21.1884945678535, 20.7287656384094, 20.5519701720443, 
    21.5739905222116, 21.8918679417571,
  18.9303526457191, 20.274712232161, 18.5138636658047, 19.7395569607073, 
    24.0947493074038, 27.0132083681126, 20.0226633238028, 20.1367588990632, 
    22.7872034912004, 20.7210183849924,
  20.4901898046254, 19.4469634862646, 21.1837070417692, 22.2330715581752, 
    21.8094416022961, 21.826933616742, 20.3538456552621, 23.8340934109302, 
    22.4198664982303, 23.159836327862,
  19.9109999486901, 23.1146421700718, 21.069002697698, 22.7342084556763, 
    25.9485804255021, 25.7840724811683, 21.5779668002319, 21.6733304774585, 
    23.4448098960645, 22.6437389538628,
  18.8270440719368, 21.5209347902249, 19.9904580994508, 20.0317053930991, 
    22.7397740352386, 25.2152921620072, 20.3247965551745, 20.1445738282327, 
    22.6303230311704, 21.4723992927257,
  22.7577045212295, 22.8924836198714, 20.3765512436531, 19.7265580707905, 
    23.9462722923718, 23.6780897041084, 20.7929154213068, 24.7557530384459, 
    22.5591589157831, 21.1946054344795,
  21.5855194202003, 20.2291006025195, 20.1297525971776, 20.3210070749892, 
    25.6053189508697, 23.1723017042731, 19.0047680771155, 17.4435336214775, 
    22.1520591139627, 20.7037993986189,
  22.7515313482526, 23.2084007855257, 22.4721595899773, 21.1291219453809, 
    24.3775544884761, 24.0538200711355, 23.5831955092598, 25.4347582314583, 
    23.3588427864257, 20.9169930185815,
  23.7907055856335, 19.4519354717177, 19.4783769827082, 22.4612060958189, 
    27.5748251455028, 25.4824865719166, 21.4506273693519, 19.2100090384522, 
    19.89619512539, 23.299806642344,
  25.111891927803, 21.5132837197623, 21.7500097380285, 20.6060950351156, 
    28.4753945980444, 24.6068237437669, 21.7917345077839, 22.4691531588236, 
    22.6220126882895, 25.3318696231738,
  20.7442210355058, 20.9202479783407, 21.1153789658916, 17.9207896412762, 
    25.1659119350521, 20.9875455685764, 22.1249484381985, 21.2292954318962, 
    22.2663908996063, 21.7409494037806,
  23.1205489231407, 19.2676046243686, 17.5607710161048, 23.4187315437524, 
    22.9455023977206, 24.5274901945454, 22.9793825028376, 22.2073551646713, 
    21.7347185842604, 23.595101659263,
  19.1916879140118, 23.0133068540555, 21.6115419472856, 19.1933684987948, 
    23.5978976623249, 22.6964834666025, 19.5108086251053, 21.0349269595516, 
    21.7579762654277, 21.5528073061353,
  22.9277871084275, 21.9051640209088, 23.8403580838155, 20.8735063410981, 
    25.1652982193381, 27.5208010146048, 23.9095662835657, 20.6301378771404, 
    21.6853926403614, 19.9115813570846,
  19.7815818650276, 20.2578502431037, 20.5399011483495, 21.5458228334826, 
    22.9288588754644, 22.7092568694927, 17.3507266016562, 19.4994848336919, 
    21.1851347356667, 21.2399054948425,
  22.5964397423441, 21.3946704378723, 18.5309597648049, 19.3290635971545, 
    25.7438307171146, 21.9221960983837, 21.5402190712922, 22.0383802890004, 
    24.8211040962597, 21.2215289624997,
  17.5922184071813, 20.759064439412, 20.6546141009909, 19.6886307764856, 
    25.6808063187578, 23.1510535079261, 22.8712711968223, 19.3646759447285, 
    22.6689817782165, 19.9233098446201,
  20.8354643524143, 23.6361190421795, 22.4199715307098, 20.1779134724923, 
    27.0529119575152, 24.9912299342735, 20.4431221715749, 22.1093939845954, 
    25.4371346503502, 21.4228002365233,
  22.9138956784773, 20.8562383479874, 17.95074971464, 19.9736909960965, 
    21.0588960911441, 24.8208840276475, 20.1645603607664, 19.5847520450156, 
    21.0587843358757, 19.8497875725498,
  22.7818670964183, 22.3395203087639, 20.7764533387754, 23.2461173308604, 
    23.9147078575073, 24.6795004378773, 21.0709413347645, 20.0156080696363, 
    20.3450168070492, 20.1298916455193,
  23.0990408015651, 21.3808923689403, 20.7044906986339, 21.6399686332365, 
    22.9757438995281, 24.0945608414141, 19.1619498115214, 20.3509308633864, 
    21.2226719751707, 20.8107919051927,
  21.3883947264998, 18.6645226899255, 18.7726631792144, 20.6799956403615, 
    23.3869340718694, 21.326622058579, 19.5958226237815, 19.0688940594358, 
    21.3093015763965, 20.1684627735478,
  23.6832578356919, 23.053614718683, 21.1197987999292, 19.8702813778058, 
    27.7948683774733, 23.3355529064126, 20.7504517556289, 20.2041484261943, 
    23.0113418092628, 24.7563485881934,
  18.8837997055759, 20.4331894915445, 17.5182077163017, 22.496635270509, 
    25.9608175792243, 26.5377502645297, 19.9552466814189, 21.8030903144122, 
    19.0665213675885, 18.7543067718812,
  20.0250381122438, 20.1199369190811, 19.1917952382023, 21.8652623827969, 
    24.5982699501338, 25.6161856135793, 21.8629025669199, 25.6641373229567, 
    24.8618367177074, 21.4505479892448,
  20.8032959402899, 19.7887632542652, 19.6712745051671, 20.4463911383844, 
    22.5115290071888, 23.5605356089489, 22.853651019952, 21.3770438985308, 
    24.695375515175, 24.3521673940476,
  25.2419423072122, 23.3806283884698, 21.3664774119649, 21.8441988502125, 
    26.0287014725512, 25.3661220308473, 24.2142324830088, 23.3476084229793, 
    20.3730372035093, 25.4221466819232,
  21.4853826267426, 17.8054985116432, 17.9022176905336, 19.2112048069753, 
    24.0963742499947, 23.1106736410241, 18.1015670118515, 23.2491976446834, 
    23.0802988884883, 23.1123266446163,
  21.9328292171759, 21.9774810864094, 18.3679346757487, 22.0913502988411, 
    25.2470978405102, 23.4092013698959, 20.2939748215147, 21.984591683745, 
    19.9427574782358, 20.1061379470214,
  19.7626479972023, 19.3279796093286, 19.83340940422, 19.2837295899993, 
    21.976933480482, 24.2480953101215, 20.2717183125162, 18.8803865569304, 
    19.1242811008471, 20.1097455121858,
  23.8564098314084, 21.1668277858941, 20.0240831662372, 21.5418250945561, 
    22.6356530714867, 22.7141614831907, 21.6842494447522, 20.6130800926184, 
    22.6489495822645, 23.408165052098,
  20.6729865378582, 20.8537223533377, 21.1355224713282, 23.0580503183898, 
    24.6126570419189, 24.3087696028367, 21.8609226532723, 19.3738110371616, 
    20.7183392418525, 17.1943845136736,
  21.9754356299466, 24.1526505016423, 20.1335340651607, 17.969718278654, 
    25.2500850270191, 24.9541013648527, 20.4825040712412, 21.8987932320236, 
    24.063161625578, 21.0237947107695,
  20.3507973364231, 20.2876377901728, 22.0607960597752, 22.9321922655592, 
    23.6116535263327, 23.4024293343729, 23.7430982539712, 21.674057222384, 
    20.1279801770363, 22.9708330866084,
  21.7558515255225, 21.0371909755942, 20.4938345994407, 23.5469447578193, 
    23.3411897185886, 23.7160074620787, 19.6137473065506, 21.9660916763639, 
    20.2147719025996, 23.1688196917367,
  21.7281427835059, 23.2686818363886, 23.1849799655181, 21.8168365830046, 
    23.8837990435528, 23.2025970466571, 20.6928624149478, 20.4076469749171, 
    20.9224852938827, 20.9193819203914,
  21.4918799517991, 21.2301998786606, 21.9239384770299, 19.0974967448306, 
    24.3132509452142, 24.1000444790023, 21.3924108559252, 22.074913607882, 
    20.9389256157484, 18.4351476450387,
  20.9502336727033, 23.2428631399006, 19.8244847927124, 19.7314076566805, 
    24.4101600701403, 25.4865561844051, 18.743828246976, 19.9186229460501, 
    20.109581246934, 20.7637994414848,
  21.095239268298, 18.9444409010423, 20.2007975816319, 18.2232780566479, 
    20.7744509759258, 24.1641729796988, 18.070447937791, 23.8005956839037, 
    20.74171196963, 20.2793228256752,
  21.9388852114143, 22.1817722537807, 20.3136043930983, 22.4978534144964, 
    22.4673751262439, 26.6514648321599, 22.5973835810623, 23.2237935475328, 
    19.6269002471305, 22.2634203309927,
  22.2374129466093, 18.40997062846, 19.2502084693846, 23.4754832850181, 
    22.4980083381104, 24.3055113609853, 18.6973926834582, 22.3003554915436, 
    24.7807601477012, 23.1447857624952,
  23.7035729991945, 19.3311878647855, 20.508799781778, 17.3901930351232, 
    23.2572851902815, 18.8414833854692, 18.1364588321687, 21.3376262193253, 
    20.6413159267135, 19.6317846891209,
  20.8478289163151, 21.1309773542641, 20.92609021264, 20.8112487342858, 
    22.7711910465343, 26.7824171857389, 22.1817490157408, 20.5732088315114, 
    20.4348870047174, 20.5253647690031,
  21.9230279401832, 21.0288957077308, 18.2782314447954, 18.0714517137996, 
    23.8700189834806, 22.6642194102985, 19.1923687690299, 23.4957527563328, 
    24.3502677257662, 22.7112981952064,
  21.5091513509786, 20.0405441367306, 20.7422503069809, 21.4063885127634, 
    23.6072660974002, 21.4273784796727, 18.8004205675483, 18.4501294853611, 
    22.8816533388277, 22.3049409113901,
  22.8833016853282, 22.1737296620837, 19.32130848855, 19.1294750863478, 
    25.5957003390634, 28.3818061542751, 22.7806783138376, 24.5400363756961, 
    21.6247477164523, 22.7657164002058,
  23.8743217377005, 22.0114193762634, 19.7555736222735, 21.1554732098952, 
    23.6169246118331, 22.4402988504091, 25.1399473788934, 23.5325500003595, 
    22.7778991433063, 21.7662183570731,
  19.6859100391343, 20.7971689298963, 19.7083366639718, 19.0123658950741, 
    22.2529400200916, 21.7718065659624, 24.1246133513329, 19.6810366313335, 
    22.7596525274184, 21.4878123586797,
  22.1954785541166, 23.2639142545952, 18.511090695693, 20.7634091483064, 
    25.4678399658171, 25.1097369803098, 19.9757105676934, 17.3930510131201, 
    22.917278188106, 24.1223364781252,
  21.4388534546269, 18.1157805576587, 18.5709920331443, 21.6804246955495, 
    21.2139919134426, 22.546855809883, 18.9471094082578, 23.4595683017459, 
    21.5302331572382, 21.3501078114966,
  17.26683273414, 21.1370727063678, 19.3753620516732, 19.046239909969, 
    23.1662841626736, 21.1900312639175, 17.8102819953445, 20.7499469089172, 
    21.6047775154296, 17.6823163689093,
  23.3476739592285, 19.8707648220565, 19.0656046238931, 20.796154385968, 
    23.1113475817135, 24.089223303911, 21.2864646471007, 20.3840094416579, 
    21.8008781868028, 25.3540031769062,
  21.2881624371116, 22.0122107198562, 21.730311044844, 17.8377915917329, 
    27.3778341561663, 24.2858122793384, 22.6159533843165, 19.2211187788598, 
    22.4040644780388, 21.9266555278908,
  23.3039946704323, 22.2387894071931, 22.8586967179414, 22.0820037773226, 
    21.5565464727976, 21.7182457145464, 23.0991458394485, 23.3873403385416, 
    21.1765921861736, 21.2394105845464,
  19.1031051229743, 19.5683892027788, 15.4653265529215, 18.9074890098494, 
    21.768261061126, 24.3881046843057, 19.1950166046849, 20.3055183675387, 
    19.534395780303, 19.2947637240416,
  21.5127971956888, 19.0942069292715, 19.3767338251079, 19.9314398111805, 
    22.1936038580888, 19.8826550781544, 18.1020532826583, 19.8294469220733, 
    21.4511967687784, 21.0823240966189,
  17.9598771434618, 22.6622790912421, 19.5293293103786, 22.5520255200037, 
    23.0784073915057, 19.790196313872, 21.7677606721171, 23.2239941759227, 
    19.0590156544851, 21.4621393605564,
  22.1909746166354, 21.9727634251639, 20.6491145877208, 23.5587539366682, 
    26.5125813123843, 24.319495408068, 22.410082317428, 20.7775520334141, 
    24.4614657447189, 22.1806566293697,
  21.8892098675853, 24.3182858015591, 21.4425994038261, 21.9268170571873, 
    21.1392127053833, 23.6146116347725, 22.131995808754, 20.8514294238815, 
    21.5294006502111, 21.0116230759699,
  21.9795025034094, 22.2059301424604, 21.4164228709442, 24.0428528268146, 
    25.9278313072514, 20.7317997839585, 20.6998410165362, 20.9934479080217, 
    21.1728705830868, 22.9764843364179,
  21.7928940416981, 21.2933391329909, 17.872251172829, 21.1322692332066, 
    24.1096714257921, 22.6547942765076, 19.6404337945902, 21.9998390726573, 
    20.3284308394674, 18.5992568079703,
  19.7215765872038, 18.3850168529869, 20.0727119027137, 18.5163558107911, 
    22.7609934018589, 23.199092566963, 17.9461966842235, 20.3829728828704, 
    21.5454714727927, 22.0478721103556,
  23.9560867394975, 22.0063139312341, 21.2659405229382, 20.7850419997789, 
    28.6300101016033, 23.7952028337735, 21.6738320150245, 23.9321434167417, 
    19.9587057147127, 24.539415188482,
  20.9293250177577, 21.9854251456441, 19.5649897527594, 17.4063341713351, 
    26.127267329833, 22.606777828558, 20.5326510473124, 23.7618595225158, 
    21.8271353276463, 22.1052069281226,
  22.4819869416745, 23.3319271939814, 21.3147553897846, 20.3313275831611, 
    25.6753800045529, 23.7378322073609, 19.2357315613588, 24.4222449595183, 
    23.4946135301726, 21.0267498828187,
  22.7426943587826, 21.9754515041939, 20.6509056465647, 21.0441984510562, 
    24.9134737010338, 25.6472424351966, 22.6718983785015, 23.4101123160913, 
    25.8606869788004, 20.8909353883345,
  21.0258747198133, 21.6175729785806, 20.1710217661128, 21.2819290142989, 
    23.2267957607011, 24.5383052359175, 21.4248017915207, 19.5733660539257, 
    22.5248211359096, 22.9996005700087,
  22.5695496548817, 21.2923015109917, 19.8556821363221, 20.2849221101071, 
    25.6669865798249, 24.062872671881, 21.3016953275113, 23.942420384798, 
    23.3974916098512, 20.5374022320011,
  23.2637821061396, 20.7527927947456, 20.2141019062476, 20.0657629076572, 
    24.6813931042881, 25.3282426359107, 19.4181731679441, 19.041336255628, 
    22.2662257916345, 23.455035383773,
  18.3830568792931, 19.6233534480576, 19.9052050179246, 19.0885324141285, 
    23.634925025883, 23.6980571037089, 19.4220461913667, 18.2622993323682, 
    22.0097588165459, 19.0971642926965,
  21.0108737753371, 21.062285221296, 18.8090368459474, 19.879499110917, 
    23.3657626307978, 22.9856512745162, 22.8544282466823, 20.9522510562678, 
    24.2189866221385, 25.0519561316447,
  21.3383089184317, 21.0799039620723, 21.6905754143959, 22.6046387078865, 
    25.1886902734136, 29.3868579563218, 23.2324725367357, 22.273800540138, 
    22.4404346740774, 21.4606606250737,
  19.1228663335468, 21.3628985966528, 20.3789071887151, 19.2116996482182, 
    24.4232718576629, 24.3804768964593, 22.6082008214178, 19.8056876628566, 
    21.7538607110906, 21.9447908762497,
  21.7443621592944, 22.9018293462479, 22.1482769972526, 22.1899843243323, 
    27.0902213163752, 25.4097675374233, 21.5907775478126, 21.6342836995343, 
    24.1180307305221, 23.7254818058622,
  19.5487232023931, 20.7029803535127, 22.2758835459625, 20.111149595995, 
    27.1193706845175, 23.9059287639524, 21.9127916090235, 20.9499683333024, 
    21.9775492639704, 21.8804881567001 ;

 concentration_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mean_source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_phase_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wind_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 concentration_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 mean_source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_phase_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 wind_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 location = 0, 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9 ;

 time = 41.666666666666667 ;

 advance_to_time = 41.666666666666667 ;
}
