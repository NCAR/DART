netcdf sgp30smosE13.b1 {
dimensions:
	time = UNLIMITED ; // (3696 currently)
variables:
	int base_time ;
		base_time:string = "1-May-2003,0:00:00 GMT" ;
		base_time:long_name = "Base time in Epoch" ;
		base_time:units = "seconds since 1970-1-1 0:00:00 0:00" ;
	double time_offset(time) ;
		time_offset:long_name = "Time offset from base_time" ;
		time_offset:units = "seconds since 2003-05-01 00:00:00 0:00" ;
	float wspd(time) ;
		wspd:long_name = "Wind Speed" ;
		wspd:units = "m/s" ;
		wspd:valid_min = 0.f ;
		wspd:valid_max = 45.f ;
		wspd:resolution = 0.01f ;
		wspd:missing_value = -9999.f ;
		wspd:threshold = "1.00 m/s" ;
		wspd:uncertainty = "+/- 1% for 2.5 to 30 m/s\n",
    "- 0.12 to +0.02 m/s at 2.0 m/s\n",
    "- 0.22 to +0.00 m/s at 1.5 m/s\n",
    "- 0.31 to -0.20 m/s at 1.0 m/s\n",
    "- 0.51 to -0.49 m/s at 0.5 m/s\n",
    "Error included in uncertainty are calibration accuracy,\n",
    "data logger timebase accuracy, and bias by underestimation\n",
    "due to threshold.  The latter assumes normal distibution\n",
    "of winds about the mean with standard deviations ranging\n",
    "between 0.25 and 1.00 m/s." ;
	int qc_wspd(time) ;
		qc_wspd:long_name = "Quality check results on field: Wind Speed" ;
		qc_wspd:units = "unitless" ;
	float wspd_va(time) ;
		wspd_va:long_name = "Wind Speed (vector averaged)" ;
		wspd_va:units = "m/s" ;
		wspd_va:valid_min = 0.f ;
		wspd_va:valid_max = 45.f ;
		wspd_va:resolution = 0.01f ;
		wspd_va:missing_value = -9999.f ;
	int qc_wspd_va(time) ;
		qc_wspd_va:long_name = "Quality check results on field: Wind Speed (vector averaged)" ;
		qc_wspd_va:units = "unitless" ;
	float wdir(time) ;
		wdir:long_name = "Wind Direction" ;
		wdir:units = "deg" ;
		wdir:valid_min = 0.f ;
		wdir:valid_max = 360.f ;
		wdir:resolution = 0.1f ;
		wdir:missing_value = -9999.f ;
		wdir:threshold = "Wind speed </= 1.00 m/s" ;
		wdir:uncertainty = "+/- 5.0 deg for wind speed > 1.0 m/s\n",
    "+/- 180.0 deg for wind speed </= 1.0 m/s\n",
    "Errors included in uncertainty are sensor accuracy,\n",
    "alignment accuracy, and A/D conversion accuracy." ;
	int qc_wdir(time) ;
		qc_wdir:long_name = "Quality check results on field: Wind Direction" ;
		qc_wdir:units = "unitless" ;
	float sd_deg(time) ;
		sd_deg:long_name = "Standard Deviation of wind direction" ;
		sd_deg:units = "deg" ;
		sd_deg:valid_min = 0.f ;
		sd_deg:valid_max = 90.f ;
		sd_deg:resolution = 0.1f ;
		sd_deg:missing_value = -9999.f ;
	int qc_sd_deg(time) ;
		qc_sd_deg:long_name = "Quality check results on field: Standard Deviation of wind direction" ;
		qc_sd_deg:units = "unitless" ;
	float temp(time) ;
		temp:long_name = "Temperature" ;
		temp:units = "C" ;
		temp:valid_min = -40.f ;
		temp:valid_max = 50.f ;
		temp:resolution = 0.01f ;
		temp:missing_value = -9999.f ;
		temp:uncertainty = "+/- 0.45 C for wind speed >/= 6.00 m/s\n",
    "+/- 0.89 C for wind speed = 3.00 m/s\n",
    "+/- 1.46 C for wind speed = 2.00 m/s\n",
    "+/- 3.07 C for wind speed = 1.00 m/s\n",
    "Errors included in uncertainty are radiation error, sensor\n",
    "interchangeability, bridge resistor precision, and polynomial\n",
    "curve fitting.  Radiation error is the largest contributor to\n",
    "the latter uncertainties.  Future algorithm development may\n",
    "reduce these uncertainties." ;
	int qc_temp(time) ;
		qc_temp:long_name = "Quality check results on field: Temperature" ;
		qc_temp:units = "unitless" ;
	float rh(time) ;
		rh:long_name = "Relative Humidity" ;
		rh:units = "%" ;
		rh:valid_min = -2.f ;
		rh:valid_max = 104.f ;
		rh:resolution = 0.1f ;
		rh:missing_value = -9999.f ;
		rh:uncertainty = "+/- 2.06 % RH for 0 to 90 % RH\n",
    "+/- 3.04 % RH for 90 to 100 % RH\n",
    "Errors included in uncertainty are calibration uncertainty,\n",
    "repeatability, temperature dependence, long term (1 yr)\n",
    "stability, and A/D conversion accuracy.  Wind speed dependence\n",
    "and radiation dependence have not been considered and may\n",
    "increase the uncertainty." ;
	int qc_rh(time) ;
		qc_rh:long_name = "Quality check results on field: Relative Humidity" ;
		qc_rh:units = "unitless" ;
	float vap_pres(time) ;
		vap_pres:long_name = "Vapor Pressure" ;
		vap_pres:units = "kPa" ;
		vap_pres:valid_min = 0.f ;
		vap_pres:valid_max = 10.f ;
		vap_pres:resolution = 0.001f ;
		vap_pres:missing_value = -9999.f ;
	int qc_vap_pres(time) ;
		qc_vap_pres:long_name = "Quality check results on field: Vapor Pressure" ;
		qc_vap_pres:units = "unitless" ;
	float bar_pres(time) ;
		bar_pres:long_name = "Barometric Pressure" ;
		bar_pres:units = "kPa" ;
		bar_pres:valid_min = 80.f ;
		bar_pres:valid_max = 110.f ;
		bar_pres:resolution = 0.01f ;
		bar_pres:missing_value = -9999.f ;
		bar_pres:uncertainty = "+/- 0.035 kPa\n",
    "Errors included in uncertainty are linearity, hysteresis,\n",
    "repeatability, calibration uncertainty, temperature dependence,\n",
    "and long-term (1 yr) stability.  Wind speed dependence has not\n",
    "been considered and may increase the uncertainty." ;
	int qc_bar_pres(time) ;
		qc_bar_pres:long_name = "Quality check results on field: Barometric Pressure" ;
		qc_bar_pres:units = "unitless" ;
	float snow(time) ;
		snow:long_name = "Snow Depth" ;
		snow:units = "mm" ;
		snow:valid_min = -25.f ;
		snow:valid_max = 1500.f ;
		snow:resolution = 0.1f ;
		snow:missing_value = -9999.f ;
		snow:uncertainty = "+/- 10.0 mm plus any offset error\n",
    "(Specified accuracy)" ;
	int qc_snow(time) ;
		qc_snow:long_name = "Quality check results on field: Snow Depth" ;
		qc_snow:units = "unitless" ;
	float snow_sen(time) ;
		snow_sen:long_name = "Snow Depth Sensor" ;
		snow_sen:units = "on/off" ;
		snow_sen:valid_min = 0.f ;
		snow_sen:valid_max = 1.f ;
		snow_sen:missing_value = -9999.f ;
	int qc_snow_sen(time) ;
		qc_snow_sen:long_name = "Quality check results on field: Snow Depth Sensor" ;
		qc_snow_sen:units = "unitless" ;
	float precip(time) ;
		precip:long_name = "Precipitation Total" ;
		precip:units = "mm" ;
		precip:valid_min = 0.f ;
		precip:valid_max = 150.f ;
		precip:resolution = 0.001f ;
		precip:missing_value = -9999.f ;
		precip:uncertainty = "Under normal conditions, uncertainty for\n",
    "rain is +/- 0.254 mm (one bucket).  Uncertainty increases to\n",
    "an unknown value during strong winds or very heavy rains (in\n",
    "excess of 75 mm per hour). The instrument is not considered\n",
    "reliable for snow amounts." ;
	int qc_precip(time) ;
		qc_precip:long_name = "Quality check results on field: Precipitation Total" ;
		qc_precip:units = "unitless" ;
	float vbat(time) ;
		vbat:long_name = "Battery Voltage" ;
		vbat:units = "V" ;
		vbat:valid_min = 9.6f ;
		vbat:valid_max = 16.f ;
		vbat:resolution = 0.01f ;
		vbat:missing_value = -9999.f ;
		vbat:comment = "This is the voltage of the CR10X battery for QA/QC purposes" ;
	int qc_vbat(time) ;
		qc_vbat:long_name = "Quality check results on field: Battery Voltage" ;
		qc_vbat:units = "unitless" ;
	float sd_wspd(time) ;
		sd_wspd:long_name = "Standard Deviation of Wind Speed" ;
		sd_wspd:units = "m/s" ;
		sd_wspd:valid_min = 0.f ;
		sd_wspd:valid_max = 9.f ;
		sd_wspd:resolution = 0.01f ;
		sd_wspd:missing_value = -9999.f ;
	int qc_sd_wspd(time) ;
		qc_sd_wspd:long_name = "Quality check results on field: Standard Deviation of Wind Speed" ;
		qc_sd_wspd:units = "unitless" ;
	float sd_temp(time) ;
		sd_temp:long_name = "Standard Deviation of Temperature" ;
		sd_temp:units = "C" ;
		sd_temp:valid_min = 0.f ;
		sd_temp:valid_max = 2.f ;
		sd_temp:resolution = 0.01f ;
		sd_temp:missing_value = -9999.f ;
	int qc_sd_temp(time) ;
		qc_sd_temp:long_name = "Quality check results on field: Standard Deviation of Temperature" ;
		qc_sd_temp:units = "unitless" ;
	float sd_rh(time) ;
		sd_rh:long_name = "Standard Deviation of Relative Humidity" ;
		sd_rh:units = "%" ;
		sd_rh:valid_min = 0.f ;
		sd_rh:valid_max = 20.f ;
		sd_rh:resolution = 0.1f ;
		sd_rh:missing_value = -9999.f ;
	int qc_sd_rh(time) ;
		qc_sd_rh:long_name = "Quality check results on field: Standard Deviation of Relative Humidity" ;
		qc_sd_rh:units = "unitless" ;
	float sd_vap_pres(time) ;
		sd_vap_pres:long_name = "Standard Deviation of Vapor Pressure" ;
		sd_vap_pres:units = "kPa" ;
		sd_vap_pres:valid_min = 0.f ;
		sd_vap_pres:resolution = 0.001f ;
		sd_vap_pres:missing_value = -9999.f ;
	int qc_sd_vap_pres(time) ;
		qc_sd_vap_pres:long_name = "Quality check results on field: Standard Deviation of Vapor Pressure" ;
		qc_sd_vap_pres:units = "unitless" ;
	float sd_bar_pres(time) ;
		sd_bar_pres:long_name = "Standard Deviation of Barometric Pressure" ;
		sd_bar_pres:units = "kPa" ;
		sd_bar_pres:valid_min = 0.f ;
		sd_bar_pres:resolution = 0.01f ;
		sd_bar_pres:missing_value = -9999.f ;
	int qc_sd_bar_pres(time) ;
		qc_sd_bar_pres:long_name = "Quality check results on field: Standard Deviation of Barometric Pressure" ;
		qc_sd_bar_pres:units = "unitless" ;
	float lat ;
		lat:long_name = "north latitude" ;
		lat:units = "degrees" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
	float lon ;
		lon:long_name = "east longitude" ;
		lon:units = "degrees" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
	float alt ;
		alt:long_name = "altitude" ;
		alt:units = "meters above Mean Sea Level" ;
	double time(time) ;
		time:units = "seconds since 1970/01/01 00:00:00.00" ;
		time:long_name = "UNIX time" ;

// global attributes:
		:qc_method = "Standard Mentor QC" ;
		:Mentor_QC_Field_Information = "For each qc_<field> interpret the values as follows:\n",
    "\n",
    "Basic mentor QC checks:\n",
    "=======================\n",
    "A value of  0 means that no mentor QC (missing/min/max/delta) checks failed\n",
    "A value of  1 means that the sample contained a \'missing data\' value\n",
    "A value of  2 means that the sample failed the \'minimum\' check\n",
    "A value of  4 means that the sample failed the \'maximum\' check\n",
    "A value of  8 means that the sample failed the \'delta\' check\n",
    "\n",
    "  Note that the delta computation for multi-dimensioned data \n",
    "  compares the absolute value between points in the same spatial \n",
    "  location, at the next point in time. \n",
    "\n",
    "Possible Combinations of mentor QC check results:\n",
    "=================================================\n",
    "\n",
    "A value of  3 means that the sample failed the \'missing and minimum\' checks\n",
    "A value of  5 means that the sample failed the \'missing and maximum\' checks\n",
    "A value of  7 means that the sample failed the \'missing, minimum and maximum\' checks\n",
    "A value of  9 means that the sample failed the \'missing and delta\' checks\n",
    "A value of 10 means that the sample failed the \'minimum and delta\' checks\n",
    "A value of 11 means that the sample failed the \'missing, minimum and delta\' checks\n",
    "A value of 12 means that the sample failed the \'maximum and delta\' checks\n",
    "A value of 14 means that the sample failed the \'minimum, maximum and delta\' checks\n",
    "A value of 15 means that the sample failed the \'missing, minimum, maximum and delta\' checks\n",
    "\n",
    "If the associated non-QC field does not contain any mentor-specified minimum,\n",
    "maximum or delta information, we do not generate a qc_field.\n",
    "" ;
		:mqc_software = "$Id$" ;
		:proc_level = "b1" ;
		:ingest_software = " smos_ingest.c,v 7.0 2001/02/06 03:45:53 ermold Exp $" ;
		:input_source = "a1 file generated from: smos13:/data/collection/sgp/sgpsmosE13.00/1051744020.icm" ;
		:site_id = "sgp" ;
		:facility_id = "E13 : Lamont_CF1" ;
		:sample_int = "snow - every 3 minutes when temp < 10.01 deg C.\n",
    "bar press - 1 minute\n",
    "all others 1 second" ;
		:averaging_int = "30 minutes" ;
		:serial_number = "SMOS8" ;
		:comment = "The time assigned to each data point indicates the end of any\n",
    "period of averaging of the geophysical data.\n",
    "\n",
    "Altitude is in meters above Mean Sea Level." ;
		:resolution_description = "The resolution field attributes refer to the number of significant\n",
    "digits relative to the decimal point that should be used in\n",
    "calculations.  Using fewer digits might result in greater uncertainty;\n",
    "using a larger number of digits should have no effect and thus is\n",
    "unnecessary.  However, analyses based on differences in values with\n",
    "a larger number of significant digits than indicated could lead to\n",
    "erroneous results or misleading scientific conclusions.\n",
    "\n",
    "resolution for lat= 0.001\n",
    "resolution for lon = 0.001\n",
    "resolution for alt = 1" ;
		:sensor_location = "Sensors heights (above base \"alt\"):\n",
    "  10m for winds\n",
    "  2m for temp, RH, and vap pres\n",
    "  1m for bar pres" ;
		:zeb_platform = "sgp30smosE13.b1" ;
		:history = "Tue Jan 10 11:43:06 2006: ncrcat added variable time=base_time+time_offset\n",
    "Tue Jan 10 11:43:06 2006: ncrcat sgp30smosE13.b1.20030501.000000.cdf sgp30smosE13.b1.20030502.000000.cdf sgp30smosE13.b1.20030503.000000.cdf sgp30smosE13.b1.20030504.000000.cdf sgp30smosE13.b1.20030505.000000.cdf sgp30smosE13.b1.20030506.000000.cdf sgp30smosE13.b1.20030507.000000.cdf sgp30smosE13.b1.20030508.000000.cdf sgp30smosE13.b1.20030509.000000.cdf sgp30smosE13.b1.20030510.000000.cdf sgp30smosE13.b1.20030511.000000.cdf sgp30smosE13.b1.20030512.000000.cdf sgp30smosE13.b1.20030513.000000.cdf sgp30smosE13.b1.20030514.000000.cdf sgp30smosE13.b1.20030515.000000.cdf sgp30smosE13.b1.20030516.000000.cdf sgp30smosE13.b1.20030517.000000.cdf sgp30smosE13.b1.20030518.000000.cdf sgp30smosE13.b1.20030519.000000.cdf sgp30smosE13.b1.20030520.000000.cdf sgp30smosE13.b1.20030521.000000.cdf sgp30smosE13.b1.20030522.000000.cdf sgp30smosE13.b1.20030523.000000.cdf sgp30smosE13.b1.20030524.000000.cdf sgp30smosE13.b1.20030525.000000.cdf sgp30smosE13.b1.20030526.000000.cdf sgp30smosE13.b1.20030527.000000.cdf sgp30smosE13.b1.20030528.000000.cdf sgp30smosE13.b1.20030529.000000.cdf sgp30smosE13.b1.20030530.000000.cdf sgp30smosE13.b1.20030531.000000.cdf sgp30smosE13.b1.20030601.000000.cdf sgp30smosE13.b1.20030602.000000.cdf sgp30smosE13.b1.20030603.000000.cdf sgp30smosE13.b1.20030604.000000.cdf sgp30smosE13.b1.20030605.000000.cdf sgp30smosE13.b1.20030606.000000.cdf sgp30smosE13.b1.20030607.000000.cdf sgp30smosE13.b1.20030608.000000.cdf sgp30smosE13.b1.20030609.000000.cdf sgp30smosE13.b1.20030610.000000.cdf sgp30smosE13.b1.20030611.000000.cdf sgp30smosE13.b1.20030612.000000.cdf sgp30smosE13.b1.20030613.000000.cdf sgp30smosE13.b1.20030614.000000.cdf sgp30smosE13.b1.20030615.000000.cdf sgp30smosE13.b1.20030616.000000.cdf sgp30smosE13.b1.20030617.000000.cdf sgp30smosE13.b1.20030618.000000.cdf sgp30smosE13.b1.20030619.000000.cdf sgp30smosE13.b1.20030620.000000.cdf sgp30smosE13.b1.20030621.000000.cdf sgp30smosE13.b1.20030622.000000.cdf sgp30smosE13.b1.20030623.000000.cdf sgp30smosE13.b1.20030624.000000.cdf sgp30smosE13.b1.20030625.000000.cdf sgp30smosE13.b1.20030626.000000.cdf sgp30smosE13.b1.20030627.000000.cdf sgp30smosE13.b1.20030628.000000.cdf sgp30smosE13.b1.20030629.000000.cdf sgp30smosE13.b1.20030630.000000.cdf sgp30smosE13.b1.20030701.000000.cdf sgp30smosE13.b1.20030702.000000.cdf sgp30smosE13.b1.20030703.000000.cdf sgp30smosE13.b1.20030704.000000.cdf sgp30smosE13.b1.20030705.000000.cdf sgp30smosE13.b1.20030706.000000.cdf sgp30smosE13.b1.20030707.000000.cdf sgp30smosE13.b1.20030708.000000.cdf sgp30smosE13.b1.20030709.000000.cdf sgp30smosE13.b1.20030710.000000.cdf sgp30smosE13.b1.20030711.000000.cdf sgp30smosE13.b1.20030712.000000.cdf sgp30smosE13.b1.20030713.000000.cdf sgp30smosE13.b1.20030714.000000.cdf sgp30smosE13.b1.20030715.000000.cdf sgp30smosE13.b1.20030716.000000.cdf sgp30smosE13.b1.BAMEX.nc\n",
    "created by user dsmgr on machine left at 1-May-2003,3:38:31, using $State$" ;
}
