netcdf filter_input {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 80 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;

	double state(time, member, location) ;
		state:long_name = "the ensemble of model states" ;

	double state_priorinf_mean(time, location) ;
		state_priorinf_mean:long_name = "prior inflation value" ;

	double state_priorinf_sd(time, location) ;
		state_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "days" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
		:model = "Forced_Lorenz_96" ;
		:model_forcing = 8. ;
		:model_delta_t = 0.05 ;
		:model_num_state_vars = 40 ;
		:model_time_step_days = 0 ;
		:model_time_step_seconds = 3600 ;
		:model_random_forcing_amplitude = 0.1 ;
		:model_reset_forcing = "FALSE" ;
		:history = "identical (within 64bit precision) to ASCII filter_ics r1371 (circa June 2005)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 location = 0, 0.025, 0.05, 0.075, 0.1, 0.125, 0.15, 0.175, 0.2, 0.225, 0.25, 
    0.275, 0.3, 0.325, 0.35, 0.375, 0.4, 0.425, 0.45, 0.475, 0.5, 0.525, 
    0.55, 0.575, 0.6, 0.625, 0.65, 0.675, 0.7, 0.725, 0.75, 0.775, 0.8, 
    0.825, 0.85, 0.875, 0.9, 0.925, 0.95, 0.975, 0, 0.025, 0.05, 0.075, 0.1, 
    0.125, 0.15, 0.175, 0.2, 0.225, 0.25, 0.275, 0.3, 0.325, 0.35, 0.375, 
    0.4, 0.425, 0.45, 0.475, 0.5, 0.525, 0.55, 0.575, 0.6, 0.625, 0.65, 
    0.675, 0.7, 0.725, 0.75, 0.775, 0.8, 0.825, 0.85, 0.875, 0.9, 0.925, 
    0.95, 0.975 ;

 state =
  -0.286964443128385, 5.73742492999917, 2.84100158144914, -3.86381062902532, 
    0.755619333941562, 0.0742229925047959, 7.58363778029272, 
    -0.909138247617973, -3.58461133272514, -1.10998591917048, 
    8.93727035936625, 3.60465839281058, 1.39855781197867, 4.94611813667615, 
    1.96550116584291, -1.87038670962402, 2.13042017834656, 7.76996326950253, 
    0.466746961370738, -5.42556759320385, -0.150209100385033, 
    0.968053099055995, 2.74099146413443, 3.23314001748027, 5.30274741550732, 
    4.90845816500769, -2.84795162589369, 0.192459429212781, 1.91784384067655, 
    8.28457946172817, 6.10574100299259, -2.14336859151112, 0.149552566166726, 
    0.14611216053799, 4.66668228703389, 8.50791660366655, 0.989044218031345, 
    1.17756012648463, -1.42856501369119, -1.62704232242793, 8.04841927814416, 
    8.04707324228465, 8.05000163773978, 8.04968176938118, 8.04889589732237, 
    8.05224789347988, 8.04692613581556, 8.04608813874835, 8.04308028677446, 
    8.04824953192639, 8.05202951766441, 8.05170040882911, 8.04881915805264, 
    8.04914855983654, 8.05057625992788, 8.05055697454878, 8.05229937130549, 
    8.04623441991265, 8.04867331374824, 8.04883346468938, 8.04668197258517, 
    8.04946362646323, 8.04477695946038, 8.04832437065785, 8.04538246670572, 
    8.05183771199285, 8.04657845445488, 8.05071487064569, 8.04863116553597, 
    8.05128957343755, 8.05170817485253, 8.04643940984882, 8.05259559206343, 
    8.04932396100225, 8.04967283377396, 8.05036642619084, 8.05259945445749, 
    8.04565764876613, 8.0550938769449, 8.04823413009183,
  0.0640296482585316, 5.61956092904613, 3.27987916729221, -3.76943334397717, 
    0.531449062421714, -0.188381149998102, 7.71558927471514, 
    -1.02459297704287, -3.26903400563159, -1.0929494101472, 8.83664296165835, 
    3.84458388974093, 1.34559672378315, 4.88613786157956, 1.75803181900479, 
    -1.88807540569014, 1.99147950522041, 7.9866170754004, 0.200810930531716, 
    -5.29411490660327, -0.267387491896848, 0.873886459935912, 
    2.64022501478228, 3.54035488300106, 5.80388229193251, 4.38013296735721, 
    -3.01655446454571, 0.385824033428311, 2.37068501463678, 8.1950543321183, 
    6.39269358339684, -0.900186657137454, -0.0340341986632688, 
    0.16896254962214, 4.76575088721626, 8.36940267399639, 1.1634266878639, 
    1.33086271548634, -1.36277118303136, -1.7578530921157, 8.02487105125812, 
    8.02352499499109, 8.02645340255173, 8.02613351983807, 8.0253476696111, 
    8.02869965248725, 8.02337788837546, 8.02253991411665, 8.01953204529517, 
    8.02470129629933, 8.02848131129745, 8.02815216337198, 8.02527090960688, 
    8.02560031731846, 8.0270280304047, 8.0270087276522, 8.02875114646545, 
    8.02268618084102, 8.02512507328792, 8.02528521246685, 8.02313375509397, 
    8.0259153816378, 8.02122870859101, 8.02477613614665, 8.02183422284287, 
    8.02828947999579, 8.02303021002943, 8.0271666410461, 8.02508292488151, 
    8.02774134059295, 8.02815992008719, 8.02289119337979, 8.02904733962292, 
    8.02577572832949, 8.0261245927511, 8.02681821062556, 8.02905120929578, 
    8.02210942032992, 8.03154564984205, 8.0246859037942,
  -0.466723127028063, 5.02506514507971, 3.79284765477527, -3.85723565893725, 
    0.780858326820499, 0.0786239510462059, 8.03918811119441, 
    -1.14388257415078, -3.43857420077785, -0.822442003001755, 
    8.99121768354778, 3.60384922397084, 1.57097067033538, 4.95954837635496, 
    1.69017899990086, -1.81849764117002, 2.06868681176738, 8.0019119904605, 
    -0.0763982868689135, -5.25647377004406, -0.388818616921354, 
    0.744719141610456, 2.77774472424496, 3.20651954380959, 5.14811099493083, 
    5.10259900203753, -2.72747388168974, -0.182975422776097, 
    1.55966544082946, 7.69532547707739, 7.11931000716429, -0.892767983589285, 
    -0.224289810020597, 0.0908871629836758, 4.56111902520684, 
    8.24759231422414, 1.2356358089374, 0.721460260194824, -1.9193076009422, 
    -1.43718643471654, 8.03741391213502, 8.03606786148522, 8.03899624759277, 
    8.03867636416192, 8.0378905339414, 8.04124252043853, 8.03592074844939, 
    8.03508277210156, 8.03207489852817, 8.03724417709197, 8.04102415727207, 
    8.04069504166542, 8.03781377832457, 8.0381431870058, 8.03957090190862, 
    8.03955160007313, 8.04129398970393, 8.0352290302024, 8.03766792899926, 
    8.03782809121036, 8.03567659018933, 8.03845823858912, 8.03377158810293, 
    8.03731899131402, 8.03437708219213, 8.04083235233009, 8.03557307180571, 
    8.03970950044586, 8.03762578466714, 8.04028417758868, 8.04070279124311, 
    8.0354340311526, 8.04159023215042, 8.03831860780689, 8.03866746508926, 
    8.03936104556804, 8.0415940828312, 8.03465228542169, 8.04408850972288, 
    8.03722877615404,
  -0.316119196314971, 4.5746586156231, 4.56435017133119, -3.59490237889361, 
    0.45430838166211, -0.28318393411794, 8.2771523250558, -1.63759546761762, 
    -2.87217772510376, -1.46784705796792, 8.61688576559717, 4.23109208995417, 
    1.1303643762498, 4.87834638070589, 2.12165558817975, -1.83048215314772, 
    2.08864030919391, 8.23134561802559, -0.552224729137157, 
    -4.87076281892297, -0.181045336401314, 0.659883301631051, 
    2.10771792701331, 3.23979803381708, 5.73916995234779, 4.8111141671893, 
    -2.85409103867871, 0.0995587772762071, 2.06788448748567, 
    8.19887599584209, 6.75960520511818, -1.22553218407605, 
    -0.232773356050789, 0.127700952984855, 4.73637315789195, 
    8.35793285933887, 0.889677415612461, 0.819819876739247, 
    -1.92350684115442, -1.49647000180116, 8.09428479992203, 8.09293873302829, 
    8.09586714045646, 8.09554726488441, 8.09476140707965, 8.09811339848228, 
    8.09279164042467, 8.09195365824274, 8.08894579467176, 8.09411504364641, 
    8.0978950189329, 8.09756588699463, 8.09468464383548, 8.09501403837388, 
    8.09644175169591, 8.0964224664384, 8.0981648363336, 8.09209993389332, 
    8.09453878269787, 8.0946989459109, 8.09254749166794, 8.09532912700739, 
    8.09064248762151, 8.09418988261725, 8.0912479572772, 8.09770320799701, 
    8.09244395193009, 8.09658036730827, 8.09449668001392, 8.09715503845852, 
    8.09757365604285, 8.09230492382912, 8.0984610844341, 8.09518947827727, 
    8.09553832671405, 8.09623193552968, 8.09846493431302, 8.09152315925196, 
    8.10095937273998, 8.0940996465557,
  -0.313363792779709, 5.0344057816642, 3.64815748145426, -3.88991435682438, 
    0.867352615072365, 0.103265214818319, 7.69326984870172, 
    -0.946643559372899, -3.62315185508623, -0.680416152385382, 
    8.83284411519763, 3.83691643107513, 1.71946514110562, 4.92807299667657, 
    1.26300844120546, -1.87936186232103, 1.71348403198872, 8.29726279720306, 
    0.102514620371878, -4.75494487870716, 0.0686411709263333, 
    0.398418807627996, 1.72617837628121, 3.03584311850336, 5.70422164785999, 
    4.85002267712671, -2.91612653692506, 0.120964313326947, 1.95129671250282, 
    8.20254710298724, 6.67227848742659, -1.48996155088154, 
    -0.049880237817249, 0.225129325371899, 4.9075665845841, 8.30145195527867, 
    0.850198202046259, 1.10536227978364, -1.8041781241431, -1.44798617547408, 
    8.07103039940547, 8.06968431841992, 8.07261272141302, 8.07229283894562, 
    8.07150700942503, 8.07485900450272, 8.06953720895906, 8.06869924005351, 
    8.06569137147651, 8.07086064085849, 8.07464061949264, 8.07431151161038, 
    8.0714302536055, 8.07175967010837, 8.0731873724705, 8.07316807675694, 
    8.07491046063756, 8.06884549478467, 8.0712843988023, 8.07144455080104, 
    8.06929308099164, 8.07207472174804, 8.0673880685092, 8.07093547081246, 
    8.06799357828672, 8.07444883004334, 8.0691895364577, 8.07332597609641, 
    8.07124226391513, 8.07390064490943, 8.07431925666453, 8.0690504989901, 
    8.07520671311015, 8.07193508063489, 8.07228393389831, 8.07297751426912, 
    8.07521056503634, 8.06826876461975, 8.07770498791652, 8.07084525307642,
  -0.374490195842141, 5.03766738450093, 3.78659241724487, -3.75687974972257, 
    0.615669225488812, -0.0910985621215707, 7.69899110146734, 
    -0.936109803354265, -3.28644563598887, -0.572742278358168, 
    8.88686765414177, 3.6374753388971, 1.69348686482315, 4.94822367003634, 
    1.39030981638479, -1.83189428800755, 1.79935616899793, 8.28173565193267, 
    -0.338958412530597, -4.84820927060241, -0.171966214017464, 
    0.702632550018905, 2.08772147654362, 2.97104595909794, 5.33914106418475, 
    5.17888386419218, -2.46229796109584, -0.0920164991714349, 
    1.9287948067872, 8.1791205907933, 6.14918709782115, -1.89050010229189, 
    -0.175394211406401, 0.0505488750921886, 4.69151734886179, 
    8.38399423318183, 0.952415757031849, 1.13987998768979, -1.79450594713957, 
    -1.62472201614172, 7.93188339122711, 7.93053733238943, 7.9334657361497, 
    7.93314586658083, 7.93236000616396, 7.9357120003114, 7.93039023792207, 
    7.92955225835471, 7.92654439100256, 7.93171363628256, 7.93549363337943, 
    7.93516449800723, 7.93228325114106, 7.93261265428545, 7.93404036418364, 
    7.93402107443462, 7.93576347009871, 7.92969852363132, 7.93213740329769, 
    7.9322975612456, 7.93014607999169, 7.93292773305628, 7.92824107142598, 
    7.93178848260981, 7.9288465716944, 7.93530181610818, 7.93004255447823, 
    7.93417898022605, 7.93209526956242, 7.93475366602302, 7.93517226775967, 
    7.92990352003568, 7.93605968813963, 7.93278808067209, 7.93313692863101, 
    7.93383053790876, 7.9360635619156, 7.92912177004917, 7.93855798579178, 
    7.93169824135183,
  -0.135343761518508, 5.52757728515, 3.19474611006247, -3.84539054459892, 
    0.623744063148895, -0.11047741716584, 7.77350881990401, 
    -1.03001274076503, -3.59801721660366, -0.932662322238443, 
    8.76754360971738, 3.69133040992024, 1.45681762218027, 4.8713961257583, 
    1.95970994123645, -1.95118968079572, 2.10895674245644, 7.86868205221293, 
    0.804350531676538, -5.1771987151552, -0.172355450627452, 
    0.368062490275655, 2.0043122313034, 3.40441769805326, 5.98029149888215, 
    4.35067089573839, -2.98696143346515, 0.237922475946765, 2.03318773255097, 
    8.06628608451637, 6.43487435208727, -1.90599244611555, 
    -0.204089115295648, 0.00199761846781343, 4.62174647205681, 
    8.49150620652178, 1.05213805279575, 1.23868967467324, -1.4385624988981, 
    -1.71618243222562, 8.01504876188507, 8.01370269161178, 8.01663110836438, 
    8.01631124257927, 8.01552536014383, 8.01887735774404, 8.01355559864798, 
    8.01271760837352, 8.00970976373335, 8.01487898889579, 8.01865900426976, 
    8.01832988377114, 8.01544861861945, 8.01577799195574, 8.01720572734072, 
    8.01718643760114, 8.01892884355878, 8.01286388126352, 8.01530278398872, 
    8.01546291350729, 8.01331144697813, 8.0160930776104, 8.01140641743883, 
    8.01495382047739, 8.01201191322022, 8.01846718957423, 8.01320793107423, 
    8.01734434196246, 8.01526060656062, 8.01791904298548, 8.0183376278205, 
    8.01306888101147, 8.01922501880101, 8.01595343937614, 8.01630228877671, 
    8.01699590078275, 8.01922891192046, 8.01228710573348, 8.02172336485749, 
    8.0148636148858,
  -0.221094579829891, 5.11864548987145, 3.90220302160582, -3.71704439823823, 
    0.516392991579168, -0.115603688620479, 8.18413610563201, 
    -1.86107943764224, -2.79785510793398, -1.60143498659939, 
    8.28010345891973, 4.50149065755163, 1.11351899256217, 4.73205365690695, 
    1.98435699129143, -1.88348409304433, 2.04298868042316, 7.9201927917558, 
    0.347099335833057, -5.22244290060941, -0.158185633794531, 
    0.660490668812624, 2.27936454679129, 3.14438157676457, 5.4234260494027, 
    4.87820969766074, -2.7571604702295, 0.186376520084024, 1.95878237304098, 
    8.29094567050072, 6.0378173333596, -2.41960729601449, 0.0742228554497925, 
    0.0979526520105705, 4.69215650050014, 8.48950706377778, 
    0.871471028366653, 1.18318518563389, -1.54215133366903, 
    -1.60980798081125, 8.01724786414914, 8.01590178790218, 8.01883017128503, 
    8.01851030354371, 8.0177244736957, 8.02107646368634, 8.01575468226925, 
    8.0149166951383, 8.01190883706001, 8.01707813767353, 8.02085808155441, 
    8.02052897435149, 8.01764771714456, 8.01797710971695, 8.0194048151873, 
    8.01938554581455, 8.02112789289784, 8.01506297655417, 8.01750185569768, 
    8.01766201004466, 8.01551053636225, 8.01829219273736, 8.01360555903185, 
    8.0171529373898, 8.0142110273182, 8.02066629265171, 8.01540701370278, 
    8.01954341955379, 8.01745973019208, 8.02011808972947, 8.02053670793046, 
    8.01526795588395, 8.02142417795805, 8.01815254895645, 8.01850140350709, 
    8.01919497068557, 8.02142803116824, 8.01448621848306, 8.0239224419281, 
    8.0170627108084,
  -0.127848674414122, 4.96037557748627, 4.09439325800478, -3.7169794413398, 
    0.44477073910235, -0.517903303832323, 7.90882692913155, -1.0666642206845, 
    -3.29366232980753, -1.17435549449348, 8.70775867842451, 3.97445270200405, 
    1.39579966578027, 4.88690113948616, 1.60544395196399, -1.94570221278918, 
    1.84476804195198, 8.15816570161787, 0.0580129229437128, 
    -5.08897597484007, -0.219285898750457, 0.618403191055331, 
    2.07896045336838, 2.80377354702267, 5.10279806958821, 5.38273876904601, 
    -2.6006730998193, -0.214593048983533, 1.56790666784087, 7.98107568979573, 
    6.75674352514547, -1.76134324659633, -0.160830861220145, 
    0.0655408042708093, 4.72371123130701, 8.33412581269298, 1.01756196082895, 
    1.16205673852155, -1.73123391225264, -1.67316390903631, 8.00217635921211, 
    8.00083030634998, 8.00375870374915, 8.00343882661262, 8.00265299453113, 
    8.00600496758628, 8.00068321555546, 7.99984522655359, 7.99683736119599, 
    8.00200661892935, 8.00578656909758, 8.00545744810367, 8.0025762188185, 
    8.00290561853691, 8.00433331810761, 8.00431401776672, 8.00605640995417, 
    7.99999149867948, 8.00243033519976, 8.00259052111871, 8.00043905795756, 
    8.00322070798437, 7.99853406435749, 8.00208147069635, 7.99913954732734, 
    8.00559477383682, 8.000335520884, 8.00447192621972, 8.00238825546567, 
    8.00504658680702, 8.00546522193146, 8.00019648188205, 8.00635265996501, 
    8.00308105085374, 8.00342990437183, 8.00412351821651, 8.0063565115556, 
    7.99941474576516, 8.00885092254149, 8.00199119242144,
  -0.630828803709246, 5.43627636342454, 3.24620543399505, -3.87610236979625, 
    0.792150346274184, 0.423472230886097, 7.94635492602599, 
    -1.35782264094528, -3.25914098377786, -0.870869432204774, 
    8.99927360486967, 3.72491061910057, 1.56893471527963, 4.89449883707157, 
    1.28206491611211, -1.85149217784664, 1.73711148770649, 8.12827524692038, 
    -0.0689669892852399, -5.17039485522251, -0.230526547195016, 
    0.872625705593235, 2.40003728109374, 2.90277572702622, 5.09833367246078, 
    5.26305025774686, -2.63307805508293, -0.0198624909175319, 
    1.71883527834189, 8.05208982375475, 6.53450483280949, -1.95379862696421, 
    -0.0603051712043219, 0.0536360371049657, 4.69678954993608, 
    8.43381945242182, 0.969717968972933, 1.13849513208301, -1.75923491537498, 
    -1.34990814965057, 8.01179654003812, 8.0104504850817, 8.01337886012048, 
    8.01305900885251, 8.01227316803283, 8.01562515548971, 8.01030337023539, 
    8.00946539174506, 8.00645754163167, 8.01162681908036, 8.01540678135805, 
    8.01507766965267, 8.01219640710862, 8.01252581724611, 8.01395355058162, 
    8.01393423533211, 8.01567662228518, 8.00961166232548, 8.0120505848725, 
    8.01221071991494, 8.01005923513989, 8.01284086070246, 8.0081542087943, 
    8.01170162898929, 8.00875971005587, 8.01521500839062, 8.00995572881853, 
    8.01409214197707, 8.0120084310702, 8.01466678988121, 8.01508541072394, 
    8.00981667193781, 8.01597287407387, 8.01270124366078, 8.01305010130453, 
    8.01374368276829, 8.0159767019476, 8.00903490914174, 8.01847115262574, 
    8.01161141992939,
  -0.102739808224615, 5.36722693552544, 3.45151929054408, -3.81820706497525, 
    0.626331061246132, -0.165959668936378, 7.776327948616, 
    -0.750663373496991, -3.57047313847476, -0.583486640344233, 
    8.97341507974645, 3.34565887327411, 1.57893542784484, 4.94605609073503, 
    1.96097866733201, -1.85293930436856, 2.17699552172131, 7.78775567296725, 
    0.402328921104871, -5.28606791437617, -0.186326190383866, 
    0.646281045725011, 2.33302013599902, 3.18906410804611, 5.44415111056742, 
    4.87152168019193, -2.79360708394479, 0.168598192722619, 2.06083929766131, 
    8.30984790207913, 6.45712929223049, -1.27512003512896, 0.145976632791232, 
    0.249716337395298, 4.8196840748129, 8.28210502140493, 1.06995109549034, 
    1.20050891269021, -1.58285175257689, -1.70788460005891, 8.00310585335446, 
    8.00175983090214, 8.00468821497095, 8.00436831834072, 8.0035824705998, 
    8.00693447003272, 8.00161271505026, 8.00077472169174, 7.99776684607434, 
    8.00293613308638, 8.00671608477799, 8.00638698387576, 8.00350574223111, 
    8.00383515253499, 8.00526282480516, 8.00524355913602, 8.00698592379319, 
    8.00092099396618, 8.00335985807112, 8.00352005031255, 8.00136852807276, 
    8.00415020846038, 7.99946356687223, 8.00301095696047, 8.00006904209446, 
    8.00652428373544, 8.00126500450336, 8.00540143897144, 8.00331774200577, 
    8.00597613475841, 8.00639475409729, 8.00112596997224, 8.00728219386315, 
    8.00401053951108, 8.00435941935886, 8.0050529951002, 8.00728604617737, 
    8.00034423026099, 8.00978045242444, 8.00292069842956,
  -0.13447792355715, 5.34834239930401, 3.56528365776525, -3.81543679672264, 
    0.545877200711709, -0.22235801584972, 8.05755485839057, 
    -1.33291425072055, -3.33116304030286, -1.26063940147856, 
    8.76308090506941, 4.06601976783629, 1.23230579010714, 4.8806616548632, 
    2.1730061719696, -1.75704306959193, 2.19833416096285, 8.19817288733674, 
    -0.64413799176752, -4.90725494895279, -0.292941935601144, 
    0.703793414781542, 2.44151641023126, 3.28303534880948, 5.45612312831761, 
    4.71885959043764, -2.94216112058173, 0.125298737529068, 1.69352301701882, 
    7.71393251200944, 6.75288476947773, -1.97988743352849, 
    -0.391952733727964, -0.142377881383643, 4.48493688476778, 
    8.49785966265834, 1.08459828460807, 1.17664445969585, -1.54490554210801, 
    -1.72772319108767, 8.03231753753121, 8.03097146833946, 8.03389985377435, 
    8.03357998078062, 8.03279415594098, 8.03614613836923, 8.03082435784606, 
    8.02998638028816, 8.02697851580403, 8.03214779795643, 8.03592775540174, 
    8.03559864640525, 8.03271739267862, 8.03304679937955, 8.0344744989841, 
    8.03445521559478, 8.03619757976042, 8.03013264940649, 8.03257153833491, 
    8.03273169687968, 8.03058021262119, 8.03336187787487, 8.0286752273135, 
    8.0322226173504, 8.029280711471, 8.03573596594661, 8.03047668595238, 
    8.03461310378942, 8.0325294125897, 8.03518777463694, 8.03560639371352, 
    8.03033764282708, 8.03649385379709, 8.0332222237734, 8.03357108411381, 
    8.03426465401722, 8.03649770397455, 8.02955591234899, 8.03899211069828, 
    8.03213238706942,
  -0.407461039995885, 5.10723389884467, 3.66285425286099, -3.83912531791724, 
    0.690599586699175, -0.0607133483133584, 7.90507541537903, 
    -1.13243234679259, -3.44566267374706, -0.912135367070285, 
    8.83331318922197, 3.78857814323574, 1.52631470785754, 4.92612088950498, 
    1.72955672477695, -1.82217658288662, 2.0013538674158, 8.12175321005623, 
    -0.351973380527814, -4.95986882267026, -0.22650230673072, 
    0.598259454785942, 2.15818192285569, 3.04815102810978, 5.33145218299279, 
    5.10771906438178, -2.65641601566637, -0.101469205416729, 
    1.80890480007524, 8.08076354361379, 6.67616709378731, -1.31684270861207, 
    -0.161768576493729, 0.114313347510058, 4.7561838705417, 8.28985969165761, 
    0.988585746262887, 1.07580080444967, -1.84946925176551, -1.4772411850725, 
    7.98870102619755, 7.98735497708676, 7.99028339338194, 7.98996350692336, 
    7.98917762664035, 7.99252962769335, 7.98720788484638, 7.98636989003321, 
    7.98336202793752, 7.98853126398469, 7.99231127112263, 7.9919821374067, 
    7.98910088786407, 7.98943027905435, 7.99085797890857, 7.99083871112449, 
    7.99258109642091, 7.98651617308728, 7.98895502730424, 7.98911518997003, 
    7.986963713804, 7.98974536393065, 7.98505870878594, 7.98860611167065, 
    7.98566419134383, 7.99211943607445, 7.98686018396346, 7.99099660332509, 
    7.98891289925457, 7.99157131212846, 7.99198990631295, 7.98672115749636, 
    7.99287731012517, 7.98960569585291, 7.98995455698984, 7.99064816988028, 
    7.99288118398832, 7.98593938301763, 7.99537562399504, 7.98851586954955,
  -0.381795387478427, 4.74224030725068, 4.49007007715971, -3.63382618226442, 
    0.43601341146343, -0.0915011779880494, 8.23414337675392, 
    -0.545513231103005, -3.39258452855095, 0.0649785049591008, 
    9.07761200888696, 3.08656563605001, 1.84828174936028, 5.01359672599858, 
    1.08327037664391, -1.87689668339354, 1.62784004519256, 8.1979364507278, 
    -0.443761113941476, -4.86282932882057, -0.0834104342979573, 
    0.58938066585012, 2.05087667465774, 3.18450167209602, 5.59299331163759, 
    4.62281729799677, -2.97622040029005, 0.287607119228634, 1.97526764923823, 
    8.2373583057071, 6.30120096486993, -2.14280755988702, 0.0572209262122654, 
    0.161600057998816, 4.79906463985816, 8.42930263182623, 0.756734177730635, 
    1.05891273838525, -1.78636938616866, -1.40025252459196, 8.0342871117038, 
    8.03294103766543, 8.03586944852359, 8.03554958583899, 8.03476371820428, 
    8.03811571496966, 8.03279394317233, 8.03195595304546, 8.0289481093636, 
    8.0341173389044, 8.03789735598595, 8.03756823560922, 8.03468697107826, 
    8.03501635229067, 8.03644407525889, 8.03642478988706, 8.03816719681565, 
    8.03210223026505, 8.0345411365748, 8.03470126071863, 8.03254979993898, 
    8.03533144042764, 8.03064477090561, 8.03419218299506, 8.03125028129207, 
    8.03770554211695, 8.03244627961837, 8.03658268565738, 8.03449896342704, 
    8.03715739088893, 8.0375759783458, 8.03230722504943, 8.03846338657767, 
    8.03519179094571, 8.03554063689738, 8.03623424293007, 8.03846727749008, 
    8.03152547252462, 8.04096171289701, 8.03410195804603,
  -0.332717646837012, 5.04193079619466, 3.86602971901095, -3.80188615237278, 
    0.672186813369311, -0.0490259358842658, 8.03428174607174, 
    -1.41846039308356, -3.15374519228697, -1.11414472351843, 
    8.72141801251302, 4.21546336838816, 1.51862337196613, 4.94371295106637, 
    1.51532252704856, -1.82172773375564, 1.842789607494, 8.30557512841396, 
    -0.499106870791182, -4.70395182604767, -0.0119066901188128, 
    0.614640662135806, 1.92437688599423, 3.2342463499054, 5.86418416870272, 
    4.52949445611448, -2.91574139348807, 0.392288615171745, 2.44357365730144, 
    8.52562001173757, 5.84342612384891, -1.79520367452253, 
    0.0211191746447478, 0.189993832214393, 4.88621884536443, 
    8.42723261135681, 0.743159800836104, 1.24703922339627, -1.73357469652931, 
    -1.45116671376665, 8.09345597633646, 8.09210997452702, 8.09503837464854, 
    8.09471845046741, 8.09393261611256, 8.09728457309755, 8.09196288808121, 
    8.09112487672774, 8.08811699317973, 8.09328624935689, 8.09706622221638, 
    8.09673707561802, 8.09385584885841, 8.09418525180706, 8.09561293148914, 
    8.09559365580517, 8.09733603301024, 8.09127115652057, 8.09370994141552, 
    8.09387017632199, 8.09171865682605, 8.09450034987276, 8.08981371244278, 
    8.09336110909317, 8.09041914965897, 8.09687437237278, 8.09161515539374, 
    8.09575155003411, 8.09366789501619, 8.09632622991925, 8.096744873567, 
    8.09147613027061, 8.09763229482361, 8.09436066762717, 8.09470954123277, 
    8.0954031448494, 8.09763613196304, 8.09069439416581, 8.10013054129165, 
    8.09327080959639,
  0.0388769325487257, 5.25486390257216, 3.7392142673928, -3.79364742218752, 
    0.532733563811476, -0.208124416484264, 7.82383372286435, 
    -0.741602930328962, -3.55592726341466, -0.580171509529784, 
    8.99448768597686, 3.62572060273321, 1.45378659865855, 4.89392414770854, 
    1.90375249966768, -1.81998006426046, 2.05105080238361, 8.1736242734634, 
    -0.340344107515875, -4.91898236179454, -0.127604785821748, 
    0.615340441279178, 2.17004830491787, 3.20789104171403, 5.53363824323934, 
    4.60276972977512, -3.0174868226324, 0.265694301205528, 1.76813200820202, 
    7.83993109075609, 6.53723741857558, -2.11705454807207, 
    -0.0639394038597668, -0.00411377365456113, 4.52361395593614, 
    8.43856087789061, 1.17795943968394, 1.16883361719698, -1.47122586683614, 
    -1.82937128153022, 8.01036903808076, 8.00902297170891, 8.01195135026713, 
    8.01163147938676, 8.01084565063754, 8.01419765561034, 8.00887585921003, 
    8.00803788140821, 8.0050300132494, 8.01019931723956, 8.01397925581749, 
    8.01365015638513, 8.01076889770413, 8.01109830670944, 8.01252601723644, 
    8.01250672525014, 8.01424908272844, 8.00818415280843, 8.01062304102778, 
    8.01078319219413, 8.00863171958423, 8.011413355689, 8.00672672582695, 
    8.0102741167294, 8.00733220181253, 8.01378748616677, 8.0085281904058, 
    8.01266461100684, 8.01058091045273, 8.01323926826768, 8.01365789515993, 
    8.00838914066467, 8.01454536740947, 8.01127372915663, 8.01162258530885, 
    8.01231615742529, 8.01454920272631, 8.00760738601532, 8.01704363479742, 
    8.01018389618941,
  -0.223861065103591, 5.5244703245249, 3.27871102341652, -3.86532643187863, 
    0.641119724498433, -0.0611063226209302, 7.92439103054256, 
    -1.00642776694058, -3.55629760991401, -0.887591634211486, 
    8.95138030750248, 3.47966983809488, 1.35032596166453, 4.88774451706684, 
    2.26918466726258, -1.86280326729815, 2.2605021064074, 7.8900889044772, 
    0.342511308811206, -5.24042041487735, -0.158513618631176, 
    0.616863963761075, 2.17609241502981, 3.09820873242375, 5.47153341586595, 
    4.96323577411841, -2.8184634675007, 0.0828240664873134, 1.88102666487054, 
    8.1293521595938, 6.44923015381679, -1.69520904872821, 
    -0.0680345433009471, 0.0379813927705293, 4.59534567719278, 
    8.49668848651387, 1.10382672192893, 1.12746151558482, -1.53980590030219, 
    -1.71800486553545, 8.07104705031463, 8.0697009849861, 8.07262936902617, 
    8.0723095059769, 8.07152366449865, 8.07487565862735, 8.06955387395475, 
    8.06871588755992, 8.0657080347228, 8.07087731258942, 8.07465729326056, 
    8.07432818060479, 8.07144691244876, 8.07177630209675, 8.07320401461612, 
    8.07318472808853, 8.07492711247808, 8.0688621734345, 8.07130107280576, 
    8.07146120595632, 8.06930973762629, 8.07209137534729, 8.06740472886182, 
    8.07095213073487, 8.06801022690103, 8.07446549052868, 8.06920620968967, 
    8.07334261280414, 8.0712589268465, 8.07391730149796, 8.07433591474959, 
    8.06906715256652, 8.0752233675486, 8.07195173477493, 8.07230058736982, 
    8.07299417091639, 8.07522722087648, 8.06828541470468, 8.07772164953657, 
    8.0708619041021,
  -0.424419940597619, 5.16456910428301, 3.73592162707502, -3.79444193528872, 
    0.597474085785512, 0.0408580413226193, 8.01210042713691, 
    -1.3523178753161, -3.35520341364771, -1.0477793379789, 8.70376345509828, 
    3.62353986687699, 1.24774684205812, 4.79254312733434, 2.38395299884109, 
    -1.88266043959908, 2.22739528141377, 7.79030412645641, 0.62268132531925, 
    -5.24984924878282, 0.00801619356042856, 0.410458726322485, 
    1.95523256930026, 3.30256390652122, 5.84259582515959, 4.51585661588404, 
    -2.9074623381624, 0.199216553797726, 2.07518604513346, 8.10179687855279, 
    6.54621483962638, -1.37952637999239, -0.15540008541033, 0.1036394421717, 
    4.76549000016584, 8.34318330142383, 0.987599538050755, 1.13921817279372, 
    -1.81275330832328, -1.54332903840187, 8.01034072287523, 8.00899463847369, 
    8.01192304557118, 8.01160317629853, 8.01081734313434, 8.01416931522414, 
    8.00884754098644, 8.00800956100287, 8.00500170860813, 8.01017096031766, 
    8.01395095053896, 8.01362182839357, 8.01074057277349, 8.0110699673128, 
    8.01249768478089, 8.01247838001208, 8.01422078604569, 8.00815582622629, 
    8.01059473185722, 8.01075485951112, 8.00860341394117, 8.01138504676278, 
    8.00669838507295, 8.01024578761514, 8.00730389480914, 8.01375914910907, 
    8.00849988249939, 8.01263628782295, 8.01055258269086, 8.01321097021267, 
    8.01362956790352, 8.00836083727512, 8.01451700246397, 8.01124539861035, 
    8.01159425752144, 8.01228785189597, 8.01452087021604, 8.00757908352475, 
    8.01701528915812, 8.01015556299476,
  -0.155079259414083, 5.34854713421298, 3.54085631345714, -3.78738477549074, 
    0.589117099685073, -0.0807417005595954, 7.90055094660108, 
    -1.21387048132465, -3.36838506750411, -1.00124039410068, 
    8.82268986893191, 3.97827626595111, 1.53142047009208, 4.86819872887329, 
    1.32953244990774, -1.90318725643095, 1.73481781363283, 8.19915939613851, 
    -0.0400664262270537, -5.05242726501901, -0.208245892503105, 
    0.608590550456738, 2.18814887052235, 3.14402119959487, 5.49459125725193, 
    4.97085110694152, -2.81914521061979, -0.0112049953284329, 
    1.76655150729918, 8.0364226221724, 6.45835942123415, -1.96425461702627, 
    -0.19424552889526, -0.00059563584021125, 4.6042751494483, 
    8.55527081528649, 1.000805804354, 1.18583264174041, -1.45921957804876, 
    -1.67574170066907, 8.04045664380093, 8.03911061158339, 8.04203902307517, 
    8.04171912025743, 8.0409332706944, 8.04428524684869, 8.03896352484343, 
    8.03812553387399, 8.03511764664345, 8.04028689534496, 8.04406685536604, 
    8.04373772214816, 8.04085649595791, 8.04118590668815, 8.04261360031323, 
    8.04259431334888, 8.04433669224341, 8.03827180705343, 8.04071058998282, 
    8.04087082199098, 8.03871933719001, 8.04150100198931, 8.03681435335096, 
    8.0403617593708, 8.03741980839325, 8.04387502843402, 8.03861580704877, 
    8.04275222130383, 8.04066855180005, 8.04332687201916, 8.04374551618834, 
    8.0384767827876, 8.04463293816736, 8.04136133243865, 8.04171018806518, 
    8.04240380704884, 8.04463678241903, 8.03769503376067, 8.0471312077124, 
    8.04027148952802,
  -0.419327851750654, 5.09121791528085, 3.60047460458456, -3.84928848925343, 
    0.881915223998541, 0.249507693601688, 7.76840041853736, 
    -1.31541599925301, -3.30901032569679, -1.17462327618133, 
    8.68313651160969, 3.84445695336349, 1.24872299151476, 4.83182531284091, 
    2.29223792959193, -1.82778171370283, 2.2719999490175, 7.83107672136147, 
    0.529531817857335, -5.42913232130671, -0.228293267575657, 
    0.902311902434011, 2.58845541212004, 3.13046063701052, 5.3396754375346, 
    4.8990526177709, -2.92073719206588, 0.183929002033492, 1.71501979331491, 
    7.83629718629903, 6.67786911261599, -2.18775690652838, 
    -0.118449735292011, 0.0958587953123032, 4.79808929133653, 
    8.34927154495326, 0.80364219920212, 1.12861356686616, -1.79399764916516, 
    -1.34074593627262, 8.04986150557355, 8.04851544705171, 8.05144386117826, 
    8.05112397532043, 8.05033810421395, 8.05369010583979, 8.04836836286702, 
    8.04753037141939, 8.04452250477888, 8.04969174673355, 8.05347174738368, 
    8.05314261136091, 8.05026136491928, 8.0505907603772, 8.05201846999442, 
    8.05199920271324, 8.05374157209286, 8.04767663765168, 8.0501154994395, 
    8.05027567169861, 8.04812417480018, 8.05090583773078, 8.04621918986209, 
    8.04976658410525, 8.04682466337539, 8.05327992155409, 8.04802066926497, 
    8.05215709429322, 8.05007336606698, 8.05273178048608, 8.05315038095233, 
    8.04788163417397, 8.05403779436985, 8.05076618758675, 8.05111503657382, 
    8.05180863560109, 8.05404166780214, 8.04709986351591, 8.05653610241316, 
    8.04967635336673,
  -0.208497866324318, 5.36195712882072, 3.42761635225899, -3.81969002089249, 
    0.710744014751226, -0.0908870999736627, 7.68378987639848, 
    -1.14720757361415, -3.41714507992721, -1.2825818891772, 8.70529267313545, 
    4.01909486739806, 1.4076533111135, 4.89647604271886, 1.66594383237293, 
    -1.89429923672971, 1.96373241249185, 8.0114860332315, 0.0992775283459772, 
    -5.17873522539628, -0.286136778716296, 0.5803608236812, 2.28913949377362, 
    3.12076648124537, 5.38537319354295, 5.08220395189805, -2.71616114384803, 
    -0.0383572085449966, 1.77380952351768, 8.16662660700764, 6.2346614920585, 
    -2.16380677333348, -0.0243205973468339, 0.0711662449367179, 
    4.63764958085106, 8.53464232435143, 0.999839811511039, 1.13049844575753, 
    -1.50602510896018, -1.64329734541272, 8.04665862352278, 8.04531256470531, 
    8.04824095240119, 8.04792108433839, 8.04713523805304, 8.0504872379207, 
    8.04516545322076, 8.04432748025733, 8.04131961182772, 8.04648888156296, 
    8.05026886367301, 8.04993974909863, 8.04705848606904, 8.04738789224242, 
    8.04881560816549, 8.04879631467535, 8.05053870105167, 8.04447374495527, 
    8.04691264245715, 8.04707279566306, 8.04492130527702, 8.04770295010741, 
    8.04301629415824, 8.04656370306985, 8.04362179824209, 8.05007706333659, 
    8.04481777983668, 8.04895421008101, 8.04687048943011, 8.04952889217639, 
    8.0499474983831, 8.04467874003487, 8.0508349350677, 8.04756331514279, 
    8.04791216873108, 8.04860575503683, 8.05083879716962, 8.04389698454787, 
    8.05333322748997, 8.04647348409446,
  -0.238483502859422, 5.63057569620397, 3.1933364406075, -3.78039570782905, 
    0.499740328433402, -0.0634595749201261, 8.10214539340856, 
    -1.27403873992232, -3.32444343537605, -0.801406327012243, 
    8.86504375597161, 3.73833870318767, 1.59443110409589, 4.89834272124513, 
    1.55792159624003, -1.86049740683282, 1.92347281777012, 7.92343352743695, 
    0.0862874051490879, -5.28616184205196, -0.0903344066758661, 
    0.854334721026399, 2.45083007472785, 3.19147557385083, 5.38746264813888, 
    4.83657588028833, -2.75806978046405, 0.23777041528938, 2.04770817031979, 
    8.26271196639469, 6.26717520513363, -1.70555285499731, 0.137116403661237, 
    0.130497908508965, 4.65885104893654, 8.4326520820692, 1.18229099897655, 
    1.23694075091156, -1.46345270659091, -1.73880830694968, 7.98520139305276, 
    7.98385532763079, 7.98678373108385, 7.98646386064516, 7.98567799219464, 
    7.9890299942537, 7.98370822351815, 7.98287023256562, 7.97986237703993, 
    7.98503162979661, 7.98881162278792, 7.98848250922101, 7.98560124797716, 
    7.98593063614684, 7.98735834461685, 7.98733906892823, 7.98908145618419, 
    7.98301651741211, 7.98545539993755, 7.98561555075559, 7.98346407650152, 
    7.98624572790957, 7.98155906655047, 7.98510647025652, 7.98216456042619, 
    7.98861980847689, 7.98336054255231, 7.98749696139785, 7.98541326169929, 
    7.98807165117146, 7.98849025613666, 7.98322149566748, 7.98937768005263, 
    7.98610607131007, 7.98645491923029, 7.98714851778109, 7.98938155961576, 
    7.98243975559079, 7.99187598728535, 7.98501624588626,
  -0.384038427802128, 4.87400359212877, 4.13112601235092, -3.74435663311066, 
    0.63624060388592, -0.127067464322961, 8.10980504205815, -1.5313458777737, 
    -3.03335699283905, -1.32031403022754, 8.58471524657531, 4.08268066712864, 
    1.3286376984562, 4.87931205813121, 1.87459372901234, -1.98860189386369, 
    1.98014323120209, 8.02821744690788, 0.684226165741447, -5.15542686933704, 
    -0.0796254374258786, 0.582777114032375, 1.90588540480968, 
    3.13809685150558, 5.91602924100888, 4.51633861724175, -3.10901414445493, 
    0.402727636260083, 2.14601547762929, 8.28170867931864, 6.12624482606027, 
    -2.38447237424904, 0.0307284996257047, 0.16804140794655, 
    4.81795844618389, 8.54261832926263, 0.62377865028743, 1.06404221790631, 
    -1.68326284304626, -1.53232886048471, 8.09854063617856, 8.09719458296018, 
    8.10012297248711, 8.09980310182865, 8.09901725068134, 8.10236924588812, 
    8.09704747180286, 8.09620948895365, 8.0932016200523, 8.09837090554269, 
    8.10215084437092, 8.10182173769994, 8.09894049690416, 8.09926990892866, 
    8.10069760467119, 8.10067832164902, 8.10242068597691, 8.09635576521779, 
    8.09879462570923, 8.09895480484611, 8.09680333043483, 8.09958497911476, 
    8.09489832666271, 8.09844572841727, 8.09550380877912, 8.10195905413761, 
    8.09669978684646, 8.1008362162981, 8.09875252921318, 8.10141087454204, 
    8.10182949824933, 8.09656074698009, 8.10271695374996, 8.09944532136362, 
    8.09979418625786, 8.10048777363632, 8.10272079777924, 8.09577899726801, 
    8.10521521639074, 8.098355494905,
  -0.166068045874098, 5.13862780327941, 3.8751704930702, -3.72878503298959, 
    0.490329914230456, -0.18645606568632, 8.17117099005183, 
    -1.65442255186901, -3.22333794142916, -1.53552478243535, 
    8.38008914867366, 4.44742569673221, 1.14632747039493, 4.73571563269893, 
    1.99599901353062, -1.79192697716005, 2.09906405990151, 7.95925439847059, 
    -0.172340714949335, -5.2357163578484, -0.259123194143074, 
    0.765479635669505, 2.54531371826308, 3.21762595963087, 5.33996209762923, 
    4.96128106911, -2.77629447676058, 0.0833008048380817, 1.86971545812894, 
    8.23751195000783, 6.19221557281705, -2.1177997457761, 
    -0.00276228838178384, 0.0664044330391792, 4.67191197458283, 
    8.49438974763282, 0.955283119069574, 1.22364055143979, -1.53908586228096, 
    -1.63871153752811, 8.03963433976519, 8.03828827878922, 8.04121668996716, 
    8.04089681154579, 8.04011096280043, 8.04346293025676, 8.03814119459735, 
    8.03730320530575, 8.03429533884089, 8.03946459074822, 8.04324455254548, 
    8.04291541482366, 8.04003418506495, 8.04036359312928, 8.04179129849061, 
    8.04177200637926, 8.04351438370948, 8.03744947714856, 8.03988830663349, 
    8.04004849213742, 8.03789703531353, 8.04067867690637, 8.03599202687991, 
    8.0395394272112, 8.0365975057686, 8.04305273851201, 8.03779350743013, 
    8.0419299142242, 8.03984622978484, 8.04250456815171, 8.04292318986944, 
    8.03765447612706, 8.04381062554971, 8.04053901605626, 8.04088788214902, 
    8.04158148372099, 8.04381446981963, 8.03687270085955, 8.04630888986856, 
    8.03944918069116,
  -0.328421294209211, 5.78980139993728, 2.7690628171166, -3.81090825896437, 
    0.690858253528794, 0.18512431033226, 7.82777336301989, 
    -0.915566429714748, -3.34307260454868, -0.559215103845528, 
    9.08242743746195, 3.39277951051778, 1.53031347977803, 4.97420114748035, 
    1.82062537256818, -1.92762859623544, 2.00451949260147, 8.07080647213674, 
    -0.040769810403645, -5.08882550626881, -0.00673596494364805, 
    0.53809126644152, 2.04292911887623, 3.22383080691096, 5.66348672406028, 
    4.71014170196943, -2.94071991455615, 0.101338221484043, 1.78789327437578, 
    7.93787846424881, 6.68676443774424, -1.78040960617413, 
    -0.210094090738006, -0.0158201915590393, 4.60880041345007, 
    8.53036090453139, 1.06057092469814, 1.17515372473323, -1.49837630743336, 
    -1.56874775665732, 8.08778082709562, 8.08643474919411, 8.08936314152609, 
    8.08904328792731, 8.08825743754004, 8.09160941625007, 8.08628764845985, 
    8.08544965824891, 8.08244181816458, 8.08761107902133, 8.09139104784605, 
    8.09106193210496, 8.08818068348119, 8.08851006822486, 8.08993778044046, 
    8.08991850729479, 8.09166087182059, 8.0855959365474, 8.08803483371216, 
    8.088194977791, 8.08604350311304, 8.08882516258312, 8.08413850853731, 
    8.08768590052778, 8.08474399564956, 8.09119925282005, 8.08593999263983, 
    8.09007639174204, 8.08799269392261, 8.09065106259137, 8.0910696745045, 
    8.08580093052015, 8.09195712393404, 8.08868550604356, 8.08903436736189, 
    8.08972793991297, 8.09196098396023, 8.08501918744724, 8.09445539925249, 
    8.08759567354318,
  -0.388062628037208, 5.19751811601855, 3.65803718211491, -3.84417124014928, 
    0.784121617058671, 0.0313079029201028, 7.94925191211957, 
    -1.41438936245881, -3.20176165174772, -1.54381056933096, 8.725276925714, 
    4.3666404088449, 1.2892252356896, 4.84520860274943, 1.18910278946798, 
    -1.9309705279183, 1.52354596200875, 8.17483253710483, 
    0.00879573796764595, -4.95203836837597, 0.0510825040672072, 
    0.398098367885993, 1.86214347557891, 3.14688851343106, 5.64247904027938, 
    4.72640496734566, -2.96158100996237, 0.0655950983143755, 
    1.65907630926234, 7.80780196906477, 6.98668014280477, -1.52295987985449, 
    -0.146548600114483, 0.0642763662641792, 4.61181980385961, 
    8.41518823427294, 1.07764629517029, 0.881567549820411, -1.75000282062248, 
    -1.45469198407633, 8.09915645899519, 8.09781042163736, 8.10073880513301, 
    8.10041891697711, 8.09963307452403, 8.10298505238254, 8.09766330873046, 
    8.09682530932606, 8.09381744691283, 8.09898674462641, 8.10276667981079, 
    8.10243756440735, 8.09955632524923, 8.09988572826475, 8.10131340347383, 
    8.10129415274461, 8.10303648678712, 8.09697160339866, 8.0994104457492, 
    8.0995706323151, 8.0974191358021, 8.10020081492535, 8.09551417877172, 
    8.09906155819127, 8.09611962363399, 8.10257487345354, 8.0973156175089, 
    8.10145202098846, 8.09936836019601, 8.10202669628211, 8.10244532180746, 
    8.09717657768227, 8.10333279224333, 8.10006113198234, 8.10041002168966, 
    8.10110358399702, 8.10333662035839, 8.09639482897281, 8.10583102940524, 
    8.09897130294888,
  -0.3885679883472, 4.77294336435643, 4.03705171811863, -3.74833411822426, 
    0.863387299797618, -0.0270694972705663, 8.02101909933749, 
    -1.02640651839248, -3.4136440203805, -0.825195665705832, 
    9.09984499709827, 3.59104555532695, 1.85552067894303, 4.97547552068251, 
    0.516039280426222, -1.91031147905655, 1.31600970396433, 8.0369489850538, 
    0.204722474642665, -5.19662104344818, -0.0261427954246635, 
    0.716825033524588, 2.14919281362241, 3.12968315827265, 5.52954865312487, 
    4.82116458649386, -2.81383161029073, 0.180753747327192, 1.96386053658018, 
    8.0773395773375, 6.10708157258223, -2.0693140050482, -0.0297290475673356, 
    0.137287067960044, 4.66454398302072, 8.47439067894065, 0.912929794229752, 
    0.803240283813739, -1.83318504890117, -1.37338626579874, 
    7.97946367130637, 7.97811762567265, 7.9810460029675, 7.98072613181789, 
    7.97994028505905, 7.98329228612216, 7.9779705016171, 7.97713251747817, 
    7.97412465873084, 7.97929394801144, 7.98307390500655, 7.98274480329737, 
    7.97986354466731, 7.9801929468352, 7.98162064481722, 7.98160137185758, 
    7.9833437353412, 7.97727879981363, 7.9797176937823, 7.9798778518545, 
    7.9777263547792, 7.98050801336404, 7.9758213647489, 7.97936876612932, 
    7.97642684661355, 7.98288211269577, 7.97762282676669, 7.98175924993657, 
    7.97967555368812, 7.98233393647318, 7.98275254871505, 7.97748377980289, 
    7.9836400057561, 7.98036835903912, 7.98071722796074, 7.9814108029355, 
    7.98364385329737, 7.97670203881499, 7.98613827996205, 7.97927853161568,
  -0.224247108938625, 5.11163640228064, 3.9393217487464, -3.72868043206993, 
    0.487270708502134, -0.216727350274794, 8.23360691693549, 
    -1.57387312064244, -3.07927658192253, -1.2307088099242, 8.63824235167306, 
    4.08390934994022, 1.338247066614, 4.83425448041078, 1.92666438290137, 
    -1.86118241388842, 2.11378451089841, 7.93605312855287, 0.174002546555119, 
    -5.24297849916535, -0.242347651216374, 0.602012384514981, 
    2.32999526941258, 3.21755186758398, 5.48789521775215, 4.94167921913094, 
    -2.76105225363334, 0.0380482986994121, 1.81236341068368, 
    8.19131781336806, 6.27088963254724, -2.26540082908494, 
    0.0117256844503284, 0.0795463429575353, 4.66976566784522, 
    8.50996315727599, 0.955011470342255, 1.13874345890886, -1.59136751217085, 
    -1.69621983292949, 8.06634664916388, 8.06500056614658, 8.06792901349702, 
    8.06760913224072, 8.06682326692206, 8.07017524222011, 8.06485350698263, 
    8.06401553385725, 8.06100766902023, 8.06617684105671, 8.06995689683883, 
    8.06962772573192, 8.06674649190451, 8.0670758925916, 8.06850362960663, 
    8.06848429864984, 8.07022674741828, 8.06416177060126, 8.06660064074129, 
    8.06676078796501, 8.06460934970851, 8.06739096030259, 8.06270429395619, 
    8.06625172717722, 8.0633098215217, 8.06976506347633, 8.06450582653434, 
    8.06864224549332, 8.06655851369453, 8.06921691082117, 8.06963551149684, 
    8.06436680636997, 8.07052289385181, 8.06725132668168, 8.06760016151005, 
    8.068293811903, 8.07052676699791, 8.06358502262952, 8.07302122562414, 
    8.0661614853083,
  -0.559545835359559, 5.53499339088047, 3.00829001964562, -3.91414583878344, 
    0.819886270633062, 0.156239631442386, 7.93569181593136, 
    -1.18204735218214, -3.49676773570362, -0.969686906083521, 
    8.96178165426411, 3.8418125260518, 1.61916957916086, 4.91023782745492, 
    1.16688414651647, -1.90658408268363, 1.68529357129999, 8.11600424419713, 
    0.0229670606830839, -5.11953621568641, -0.171940107307873, 
    0.65454775070121, 2.18229064383286, 3.03808006960453, 5.37374629463594, 
    5.09607488431934, -2.73645170712769, 0.00929062581437354, 
    1.79026207594416, 8.12535745009454, 6.59444460761456, -1.71885590248065, 
    -0.00904178334794297, 0.134935980525889, 4.75546041259235, 
    8.42136555725956, 0.940640287396634, 1.09912997661105, -1.7125062138288, 
    -1.44630932638948, 8.03471240695045, 8.03336632408215, 8.03629471150327, 
    8.0359748464683, 8.03518903172979, 8.03854101561389, 8.03321922953559, 
    8.03238125279173, 8.02937338524507, 8.03454267362959, 8.03832263068523, 
    8.03799350804412, 8.03511226179597, 8.03544166696055, 8.03686937870214, 
    8.03685007651434, 8.03859245505059, 8.03252751231216, 8.03496640645098, 
    8.03512655628616, 8.03297508746723, 8.03575673583572, 8.03107009506742, 
    8.03461748692232, 8.03167559359009, 8.03813084182013, 8.03287156319871, 
    8.03700797670577, 8.03492428217655, 8.03758263605895, 8.03800125673021, 
    8.0327325124333, 8.03888872473711, 8.03561710261623, 8.0359659455038, 
    8.03665952707417, 8.03889257532727, 8.03195077616072, 8.04138697883587, 
    8.03452725119203,
  -0.30383452334819, 5.46878591446747, 3.19268278608883, -3.86077519726869, 
    0.715628067822479, 0.050594082533481, 7.71943975759205, 
    -0.904853208018582, -3.46951408555647, -0.661206589414539, 
    8.97496011587966, 3.71370016354662, 1.64355468458624, 4.95857268963752, 
    1.39141869740399, -1.8494980262044, 1.77481788955909, 8.29570612458822, 
    -0.394773493096409, -4.78323084879143, -0.0611498449021256, 
    0.494879287034204, 1.92105733108085, 3.09287071926084, 5.57625458060371, 
    5.01524056081112, -2.73947382235974, -0.100486297213065, 
    1.79897217079352, 8.09114162995688, 6.59525346365466, -1.61164581932783, 
    -0.230753627038665, 0.0389301118338327, 4.72166548794732, 
    8.4526023332752, 0.970122420174462, 1.22436619585072, -1.61194443199655, 
    -1.60601581784158, 8.01784055679242, 8.01649450622891, 8.01942288458067, 
    8.01910301523627, 8.01831717337985, 8.02166916337586, 8.01634739203725, 
    8.01550940123544, 8.01250154955667, 8.017670828647, 8.02145080509517, 
    8.02112169166515, 8.01824043082579, 8.01856981333961, 8.01999752456253, 
    8.01997824255521, 8.02172062388307, 8.0156556873019, 8.01809457615572, 
    8.01825471942745, 8.0161032398041, 8.01888487971433, 8.01419823978412, 
    8.01774564414124, 8.01480372972575, 8.02125900504165, 8.01599972296539, 
    8.02013612130195, 8.01805243215675, 8.02071080669325, 8.02112942646541, 
    8.01586066581278, 8.02201687696971, 8.01874524000816, 8.01909410477871, 
    8.01978768490431, 8.02202072320268, 8.01507891656142, 8.02451516277474, 
    8.01765540785427,
  -0.334742867549649, 5.14125461377586, 3.54230429639277, -3.77750402275756, 
    0.839453748207914, 0.1897437392207, 7.50561868519586, -1.07545435525469, 
    -3.4040046228885, -1.10390690202888, 8.66213087943711, 4.00625757816153, 
    1.40617353138252, 4.83293489530886, 1.56615075470632, -1.90189728815541, 
    1.88068318150667, 7.90284204368534, 0.171284229613737, -5.22283970601914, 
    -0.138213881939226, 0.622451386507507, 2.25664721439287, 
    3.13777989268047, 5.3944066814289, 4.99466602801937, -2.68735266403678, 
    -0.0261182161472071, 1.8623358880241, 8.11789663412045, 6.60658207544517, 
    -1.48879125489931, -0.146968874310344, 0.108390974323727, 
    4.76029322153529, 8.37780945185287, 0.983280669232855, 1.08613386226535, 
    -1.75628356163781, -1.4233047084892, 7.98303365333326, 7.98168756627967, 
    7.98461592991815, 7.98429606113214, 7.98351026353489, 7.98686226565092, 
    7.98154043919681, 7.98070245813652, 7.97769459699764, 7.98286394586738, 
    7.98664385176805, 7.98631478055322, 7.98343351607637, 7.98376293637706, 
    7.98519063024017, 7.98517135474675, 7.98691368232779, 7.9808487262477, 
    7.98328765541146, 7.98344781095829, 7.98129631188263, 7.98407798391964, 
    7.97939134576331, 7.98293872578789, 7.97999682525001, 7.98645210623096, 
    7.98119279002825, 7.98532922309045, 7.98324551868212, 7.98590385895434, 
    7.98632249203397, 7.98105371677212, 7.98721001759527, 7.98393835130047, 
    7.98428720639163, 7.98498073106078, 7.98721385056744, 7.98027200931123, 
    7.98970824455384, 7.98284852147235,
  -0.511684476546709, 5.31771817628145, 3.35829649304193, -3.84978443647909, 
    0.83914072017909, 0.257301066189067, 7.53026316547204, 
    -0.621402624289854, -3.33160255073745, -0.401536812617594, 
    9.13458892411593, 3.24214870315883, 1.64448420138002, 4.98975451910302, 
    1.37461302449055, -1.99575506426518, 1.72361822314997, 8.05265534239296, 
    0.387966705447695, -5.1321788616508, 0.071793598742365, 
    0.610020032162997, 1.94357524151375, 3.11200013038011, 5.69392869370903, 
    4.63565744106658, -2.95239469356144, 0.33623117560046, 2.10063946526153, 
    8.20470738245619, 6.4910915616897, -1.74700317278473, 
    -0.0138591897602698, 0.139893415406901, 4.81501713013068, 
    8.39395166578907, 0.959467567877372, 1.14966466423426, -1.82119631264478, 
    -1.51994466477573, 8.05120719068645, 8.04986112002189, 8.05278950073453, 
    8.05246963247795, 8.05168379597505, 8.0550357929042, 8.04971399269703, 
    8.04887600993854, 8.04586815452868, 8.05103746453144, 8.05481738612099, 
    8.05448830465927, 8.0516070421023, 8.05193644773738, 8.0533641402534, 
    8.0533448786207, 8.05508720970696, 8.04902230357999, 8.05146118300174, 
    8.0516213343784, 8.04946987549008, 8.0522515215345, 8.04756487717346, 
    8.05111225383048, 8.04817035101523, 8.05462561060981, 8.0493663239951, 
    8.05350274339931, 8.0514190539949, 8.05407742898302, 8.0544960369629, 
    8.04922728155305, 8.05538350623924, 8.0521118591405, 8.05246073976719, 
    8.05315429308545, 8.05538735036408, 8.04844551856921, 8.05788176274914, 
    8.05102204363354,
  -0.408268076442572, 5.08939247388129, 3.57015901505855, -3.88113526782714, 
    0.899105242825115, 0.151975287240508, 7.78663171238856, -1.0046374186651, 
    -3.41478645711713, -0.786681529945049, 8.92380506016963, 
    3.46089505453539, 1.50023637986822, 4.96688075239906, 2.08748334578211, 
    -1.85859733988479, 2.22345250975456, 7.90304673127716, 0.173413502291574, 
    -5.24829913013333, -0.237344986772075, 0.607022924503535, 
    2.31429802225928, 3.14433784860866, 5.39827812922273, 4.94523165580369, 
    -2.8079630670756, 0.132089336116378, 1.91091798477599, 8.33493189846732, 
    6.23863985828159, -2.07353514691034, 0.131811619386467, 
    0.242121306281741, 4.95173657178439, 8.32868186231273, 0.745910805855725, 
    1.27001047020081, -1.7947749023847, -1.40937886190185, 8.03082037934898, 
    8.02947436247971, 8.03240273314067, 8.03208287031102, 8.03129700290428, 
    8.03464900029576, 8.02932725553363, 8.02848925702118, 8.02548139165601, 
    8.03065066895091, 8.03443059517177, 8.03410148392434, 8.03122025340554, 
    8.03154964161969, 8.03297733839067, 8.0329580690656, 8.03470042664175, 
    8.02863555033528, 8.03107436872305, 8.03123457583572, 8.02908307014757, 
    8.03186474346781, 8.02717811031849, 8.03072550642043, 8.02778355262404, 
    8.03423879367774, 8.02897955246666, 8.0331159513614, 8.03103229023665, 
    8.03369062090217, 8.03410926359818, 8.02884049892219, 8.03499670037357, 
    8.03172507658764, 8.03207394180823, 8.03276754310095, 8.03500054708629, 
    8.02805875926028, 8.03749496356532, 8.03063522493568,
  -0.484227990525675, 5.13211430031823, 3.53793974163889, -3.85303467598537, 
    0.792978954351067, 0.154144728420581, 7.69971636271452, 
    -1.04814414658396, -3.38730426319906, -0.717145182053223, 
    8.83442582496264, 3.74908684751545, 1.66555034493882, 4.97902421573329, 
    1.45746989648326, -1.87073686434003, 1.80338892588112, 8.23609078664331, 
    -0.17850481773602, -4.82617343119723, 0.0530260236555174, 
    0.455142610357697, 1.94774229574462, 3.27694418358193, 5.70667097012732, 
    4.61757746485022, -2.79690815509145, 0.0601629269124873, 
    1.81501960067027, 7.86277574395838, 6.61669859127906, -1.8658974198798, 
    -0.318423401681626, -0.0215134223917905, 4.68117895351729, 
    8.40032054677791, 0.930197024640019, 1.13130494856636, -1.83630267640464, 
    -1.420500355997, 7.97758627711671, 7.97624019782646, 7.97916860666047, 
    7.978848726731, 7.97806287993768, 7.98141488178617, 7.97609310164981, 
    7.97525512889263, 7.97224725480147, 7.9774165139088, 7.98119650545008, 
    7.98086738320506, 7.97798612636129, 7.97831553155207, 7.97974325154695, 
    7.97972394750692, 7.98146634202936, 7.97540138362727, 7.97784027375253, 
    7.9780004214987, 7.97584896140629, 7.97863058637871, 7.97394393663429, 
    7.97749133789652, 7.97454943977607, 7.98100470295462, 7.97574542003841, 
    7.97988185971879, 7.97779813429999, 7.98045653006461, 7.98087513522205, 
    7.97560638877169, 7.98176256386865, 7.97849096051479, 7.97883980025854, 
    7.97953340290703, 7.98176642960928, 7.97482462679817, 7.98426086574666, 
    7.97740113282623,
  -0.254961512061245, 4.85628747772919, 4.11539982707618, -3.73795915371266, 
    0.519451038538547, -0.293205627890072, 8.01132791634584, 
    -1.10397417438693, -3.52700683416023, -0.908654435972977, 
    8.74470589724551, 3.90498886101773, 1.52679725069856, 4.87257493622702, 
    1.67972613292002, -1.85630324233558, 1.98090971128855, 8.12300480264832, 
    -0.0248989288472855, -5.05478959601003, -0.24628196373279, 
    0.489961933562502, 2.22147682166977, 3.27355308585836, 5.56749378934711, 
    4.67093214250519, -2.9271371629432, 0.11060976268921, 1.66880428437704, 
    7.72854948054199, 6.78594852837228, -2.02727605176093, 
    -0.249400551816536, 0.0248730023773532, 4.73203452733369, 
    8.37180124134064, 0.991398601329776, 1.15349481977108, -1.80727973078186, 
    -1.59406200226693, 8.00990235482796, 8.0085563067711, 8.01148470521403, 
    8.01116484521479, 8.01037896528273, 8.01373096344843, 8.00840921072705, 
    8.007571217287, 8.00456336632335, 8.00973260794477, 8.01351261390882, 
    8.01318346900384, 8.01030221953184, 8.01063161225272, 8.01205932968777, 
    8.01204005053848, 8.01378244576695, 8.00771750350474, 8.01015638728785, 
    8.01031653513492, 8.0081650450106, 8.01094669779213, 8.00626003254852, 
    8.00980745882344, 8.00686552427486, 8.01332078862845, 8.00806153838365, 
    8.01219795199627, 8.01011423839177, 8.01277263898214, 8.01319123237496, 
    8.00792249949489, 8.01407865102905, 8.01080704405099, 8.01115589305292, 
    8.01184951111934, 8.01408252745335, 8.00714072747503, 8.01657697103916, 
    8.00971721182996,
  -0.112124515138242, 4.9562688317636, 3.99821899590358, -3.78072160255053, 
    0.697930333206632, -0.209266596039841, 7.58278740538539, 
    -0.817217263462599, -3.38066582913942, -0.987021465741976, 
    8.81044736939451, 3.70070519255069, 1.38053547362605, 4.93624880531074, 
    1.94397273048135, -1.93261520002394, 2.08171040010792, 8.04838926674463, 
    0.0640099961512071, -5.11965192082412, -0.244391532119409, 
    0.424222745057574, 2.10311588543777, 3.16886778699967, 5.54340064942845, 
    5.11293428217671, -2.63810251749846, -0.204900322733424, 
    1.73132160019192, 8.17668000469939, 6.63214552962907, -2.00671694813842, 
    -0.265040230677127, 0.0372463360473547, 4.79854721180684, 
    8.48581167204031, 0.752646201873523, 1.19916976119838, -1.65976405689612, 
    -1.58659306296168, 8.05749008042156, 8.05614400514745, 8.0590724142913, 
    8.05875254901356, 8.05796668479869, 8.06131867558955, 8.05599692428337, 
    8.05515892620076, 8.05215108179316, 8.05732031859245, 8.06110032362233, 
    8.06077119242081, 8.05788993641938, 8.05821931914628, 8.05964704564377, 
    8.05962776741319, 8.06137014820016, 8.05530520154032, 8.0577440920662, 
    8.05790423167171, 8.05575275145592, 8.0585344025007, 8.05384775082814, 
    8.05739514768014, 8.05445324187867, 8.06090850968312, 8.05564926072908, 
    8.05978565882815, 8.05770193449757, 8.06036034120524, 8.06077894195633, 
    8.05551020340934, 8.06166636313573, 8.05839476278319, 8.05874360760913, 
    8.05943719795653, 8.06167023705565, 8.0547284335881, 8.06416467155828, 
    8.05730492623855,
  -0.372889120793953, 5.23296076672635, 3.59518527319873, -3.82329248498294, 
    0.683073640878727, 0.0760809057545367, 8.0429477926871, 
    -1.04278662734613, -3.33685661700594, -0.584855079993398, 
    9.01891916402909, 3.43781939368459, 1.47620188553317, 4.88087022904023, 
    1.90044435924891, -1.85809721821981, 2.07846101233416, 7.89261093849664, 
    0.304860256375378, -5.34444470548094, -0.0949210086355678, 
    0.832714995254732, 2.54485683104801, 3.34501802546281, 5.54540688439539, 
    4.79114492191789, -2.73770081281334, 0.0896837282278617, 
    1.88776560537006, 7.95784556574997, 6.65391849481067, -1.79537187041921, 
    -0.288873802970327, -0.000805357877543298, 4.69059264240158, 
    8.4177595977046, 0.950767503258712, 1.1561958876069, -1.73428807352474, 
    -1.57130793180634, 8.02433914192005, 8.02299308674288, 8.0259214823465, 
    8.02560162039352, 8.0248157563295, 8.02816775785724, 8.02284596812954, 
    8.0220079943086, 8.0190001390421, 8.02416938992553, 8.02794937638279, 
    8.02762027482672, 8.02473901178236, 8.02506842325089, 8.02649613835827, 
    8.02647683952859, 8.02821923459649, 8.02215425994566, 8.02459318125309, 
    8.02475332639492, 8.02260183858454, 8.02538347924154, 8.02069680679784, 
    8.02424422707821, 8.02130232563972, 8.02775758787755, 8.02249830656238, 
    8.02663474305841, 8.02455102754188, 8.02720941943136, 8.02762802726119, 
    8.02235925768363, 8.02851546433282, 8.02524383528119, 8.0255926930721, 
    8.02628628179363, 8.02851931735462, 8.02157752190858, 8.03101375924758, 
    8.02415401939602,
  -0.46538990884468, 5.12093201712819, 3.62491893385452, -3.86958448784451, 
    0.83298679497802, 0.0444091342105404, 7.6584705631972, -1.13580251508306, 
    -3.53090376788223, -1.39199140538999, 8.66094386417613, 3.8484759924229, 
    1.22069565425433, 4.90568842958766, 2.21761598252042, -1.95142725724117, 
    2.16063879056847, 8.08971304384538, 0.158400082964435, -5.00836670298469, 
    -0.232285238566822, 0.329330676480398, 2.02178824130958, 
    3.31302917518162, 5.73340725940784, 4.71883664611075, -2.72017024449988, 
    0.111509974683007, 2.10850116654631, 8.31458755139284, 6.21577406268846, 
    -1.80595346972883, -0.150645931490642, 0.0778432014266612, 
    4.78013018266698, 8.44974705189955, 0.755417424822593, 1.15627686987171, 
    -1.80372784312386, -1.4368271785613, 8.02555231451936, 8.02420629020087, 
    8.02713465914491, 8.02681478094748, 8.02602894531773, 8.02938093043643, 
    8.02405917252972, 8.02322118438985, 8.0202133095742, 8.02538260101025, 
    8.02916254086117, 8.02883343180498, 8.0259521908726, 8.02628160172573, 
    8.0277092873865, 8.02769000782034, 8.02943237165303, 8.02336746347433, 
    8.02580631988428, 8.02596651173347, 8.02381499733977, 8.02659667735388, 
    8.02191002817771, 8.02545742649415, 8.02251550148281, 8.0289707418063, 
    8.02371147533101, 8.02784789413191, 8.02576422130479, 8.02842256910111, 
    8.02884120289679, 8.02357243767901, 8.0297286554016, 8.02645701182523, 
    8.02680588262093, 8.02749945853186, 8.02973249494079, 8.02279070655047, 
    8.03222689582242, 8.02536716714439,
  -0.213707927849421, 4.74445521303228, 4.36243587156398, -3.56343971863069, 
    0.394713855384994, -0.132179752659896, 8.26530105703194, 
    -1.85598568118445, -3.00630823924459, -1.46573898170768, 
    8.32673988411071, 4.23095141272365, 1.06080503485006, 4.68215890725104, 
    2.361270837149, -1.83785857509418, 2.2205450876445, 7.81447005669439, 
    0.677034627973507, -5.31919432937413, -0.166993486839092, 
    0.687287769448932, 2.34065182087267, 3.14494116127578, 5.42898143290107, 
    4.95370212171025, -2.76656199199528, 0.00821863420019144, 
    1.77490221075949, 8.02113518035129, 6.73995039809122, -1.90923622967171, 
    -0.277708211745761, 0.00861597479186895, 4.71092891085868, 
    8.45268654759141, 0.8506007925405, 1.11746948031105, -1.71159225825544, 
    -1.56545498607342, 8.01534813111611, 8.01400207460825, 8.0169304727235, 
    8.01661059838674, 8.0158247270792, 8.01917673092573, 8.01385497400617, 
    8.01301697322332, 8.01000912904023, 8.01517838429971, 8.0189584098389, 
    8.01862926821463, 8.01574799913788, 8.01607737628003, 8.01750508433943, 
    8.01748583770454, 8.01922821126669, 8.01316327195821, 8.01560217078421, 
    8.01576229517988, 8.01361080249338, 8.01639247293147, 8.01170581204634, 
    8.01525321902194, 8.01231128873972, 8.01876657258601, 8.01350730550028, 
    8.01764370433029, 8.01555999064109, 8.01821842778815, 8.01863700352948, 
    8.01336825682234, 8.01952443058049, 8.01625280783506, 8.01660166361193, 
    8.01729525840292, 8.01952831785824, 8.01258649953286, 8.02202276244364, 
    8.01516297967888,
  -0.354253805253355, 5.02626213313622, 3.66369115125695, -3.8898358968592, 
    0.924303847041926, 0.14910476973298, 7.83283223981111, -1.07137368494709, 
    -3.57323331918587, -1.00613675668888, 9.01108328494785, 3.93479871514605, 
    1.56869776222918, 5.0127691334223, 1.33946690978497, -1.83863958256468, 
    1.66647698950183, 8.50652031029659, -0.366306643379336, 
    -4.53374420951913, 0.215345220798305, 0.433671646874425, 
    1.73854189264031, 3.20081133517653, 5.85055802261184, 4.7715293252243, 
    -2.84918349266145, -0.0732650723399992, 1.67757309550041, 
    7.99402180905769, 6.6234847491883, -2.26708684030716, -0.211177851608585, 
    0.0644883252850232, 4.77611082687838, 8.46830094362704, 
    0.664507166375527, 1.09547710802794, -1.68417327556992, 
    -1.43867214683855, 8.07646383959192, 8.07511777329095, 8.07804616877085, 
    8.07772630489128, 8.07694045118643, 8.08029243795847, 8.07497066556583, 
    8.07413267676143, 8.07112482570676, 8.07629409221687, 8.08007406554953, 
    8.07974495354477, 8.07686369220711, 8.07719308462944, 8.07862079480794, 
    8.07860151366932, 8.08034389568151, 8.07427896344657, 8.07671785395731, 
    8.07687799175901, 8.07472653043317, 8.07750817698691, 8.07282151394829, 
    8.07636891248975, 8.07342700279209, 8.07988226100364, 8.07462299682927, 
    8.07875940668666, 8.0766757061138, 8.0793341012917, 8.07975269517072, 
    8.07448395310798, 8.08064012505922, 8.07736851764052, 8.0777173791969, 
    8.07841097170446, 8.08064400068284, 8.07370219687075, 8.08313841796617, 
    8.0762786890214,
  -0.331880340559452, 5.5607184860511, 3.13372919810169, -3.83851932782074, 
    0.626443894247916, -0.0852939075757211, 7.72518914128875, 
    -0.969197950086559, -3.59553822315155, -1.0029722405006, 
    8.85777387931795, 3.62639626646207, 1.45720304504158, 4.90537011419966, 
    1.86106812382193, -1.89462345982372, 2.05194170403437, 7.87328950640776, 
    0.559784410297899, -5.25475351482978, -0.183412691046866, 
    0.767004113954331, 2.249826606581, 2.98651841705194, 5.33284335358057, 
    5.08867831841173, -2.69362148121182, 0.164158509551106, 2.09587743031142, 
    8.30683233413412, 6.37666892138954, -1.31042748913643, 0.117389199363156, 
    0.236351174457826, 4.84944162085223, 8.27933166282093, 1.07400921544004, 
    1.26529040655505, -1.6531327457985, -1.62742218149485, 7.98886074101116, 
    7.98751465173438, 7.99044310214058, 7.99012319948982, 7.98933734532982, 
    7.99268932028297, 7.98736760359469, 7.98652961060809, 7.98352174396273, 
    7.98869093974203, 7.99247098207231, 7.99214182188218, 7.98926058214595, 
    7.98958997188185, 7.99101768400214, 7.9909983974729, 7.99274079410412, 
    7.98667586103069, 7.98911470711471, 7.9892748692242, 7.98712340791625, 
    7.9899050608787, 7.98521841730526, 7.98876580378576, 7.98582391133563, 
    7.99227914172998, 7.98701990307211, 7.99115630975084, 7.98907259668756, 
    7.9917309901737, 7.99214960072979, 7.98688087508361, 7.99303699721681, 
    7.98976541354763, 7.99011424484412, 7.99080785783149, 7.99304087450904, 
    7.98609911509663, 7.99553530398085, 7.98867556396065,
  -0.0494056688368833, 5.5215226325288, 3.31049275092938, -3.76252882039047, 
    0.50017793401991, -0.197266996820538, 7.99052730926133, -1.0470883727397, 
    -3.42711937875077, -0.725814483554624, 8.87925969471127, 
    3.66346580454709, 1.58424593033522, 4.89985880294553, 1.6096868782791, 
    -1.8599191719451, 1.94838956838861, 8.10826808523861, 
    -0.0628669731308649, -4.98543827105502, -0.23799875592816, 
    0.45298789151246, 2.08279169391002, 3.09973113196072, 5.43124831067808, 
    5.02076554737492, -2.655872748055, -0.105840793248682, 1.77336360768584, 
    7.94570107040412, 6.69180519009989, -1.30241553844537, 
    -0.199630239399266, -0.0165862616900053, 4.49993306317681, 
    8.4131041742617, 1.24729308882402, 1.13925844855678, -1.4224815487804, 
    -1.74173448163441, 7.98213215214043, 7.98078609522424, 7.98371445883095, 
    7.98339458439711, 7.98260877595682, 7.98596076757772, 7.9806389672733, 
    7.97980099199494, 7.97679311767844, 7.98196245308289, 7.98574236478666, 
    7.98541326413493, 7.98253201582621, 7.982861443215, 7.98428913316915, 
    7.98426984840061, 7.98601218936142, 7.97994726532466, 7.98238615686924, 
    7.98254632252623, 7.98039483370167, 7.98317649174947, 7.97848985374636, 
    7.98203724355955, 7.97909533013818, 7.98555059366844, 7.98029129637848, 
    7.98442772864444, 7.98234404153511, 7.98500238518435, 7.98542100998722, 
    7.98015225858032, 7.98630850919448, 7.98303684399029, 7.98338571838762, 
    7.98407927112225, 7.98631233090106, 7.9793705121882, 7.98880673335952, 
    7.98194701182001,
  -0.444014424758751, 5.02737920833059, 3.73267594472118, -3.87361313865236, 
    0.753852067536012, -0.0158930757189786, 7.87162959922826, 
    -0.929231558928722, -3.49807382873158, -0.584452525879808, 
    8.92947758568362, 3.62022808102576, 1.66562709545661, 4.94207302211812, 
    1.55228365860228, -1.863738767573, 1.93863510487884, 8.07323793121579, 
    -0.052572227146569, -5.03064445862744, -0.128203295985514, 
    0.52770419612836, 2.0977144064392, 3.17715557666526, 5.535052200501, 
    4.64379040917751, -2.92934248815132, 0.299041949094895, 1.93915875286466, 
    8.14530354777605, 6.54789553168024, -1.94249402574132, 
    0.0963091366593622, 0.223508999493305, 4.90200580289734, 8.2724381762446, 
    0.882336803691907, 1.15617643302401, -1.90112033104901, 
    -1.49534936295466, 8.03560172444289, 8.03425572704377, 8.03718409913924, 
    8.03686421214872, 8.03607835920507, 8.03943033268555, 8.03410860490061, 
    8.03327061092619, 8.03026274015829, 8.0354320104982, 8.03921196922677, 
    8.03888284766301, 8.03600160854101, 8.03633102870606, 8.03775870836128, 
    8.03773944046976, 8.03948179978501, 8.03341689529173, 8.03585573636598, 
    8.03601594556254, 8.03386440801658, 8.03664609548498, 8.03195943699747, 
    8.03550684729393, 8.03256490613774, 8.03902014921865, 8.03376090575686, 
    8.0378973188938, 8.03581364366344, 8.03847200118023, 8.03889063214862, 
    8.0336218756123, 8.03977807504513, 8.03650641170095, 8.03685531156334, 
    8.03754887792383, 8.03978189617453, 8.03284012109511, 8.04227631297, 
    8.03541658281281,
  -0.491662054055454, 4.90673660582467, 3.93652758818775, -3.81271636586768, 
    0.754614216311681, 0.145320153220008, 7.99911886187926, 
    -1.25660017493175, -3.30606525335129, -0.833205532882565, 
    8.95831741577005, 3.78940293710389, 1.54268478236543, 4.98328591182111, 
    1.70802309404551, -1.83472321999128, 1.95694706321157, 8.24253502654278, 
    -0.447457496741195, -4.91194095166963, -0.120188956056645, 
    0.927092594009629, 2.19245837997767, 3.13462695854128, 5.65202285902552, 
    4.95695352522368, -2.62380365744065, 0.31924956135219, 2.60864370552598, 
    8.66413602141873, 5.99611911146124, -1.28857121526026, 
    -0.0230542338195771, 0.262741857344903, 5.03068440384296, 
    8.3452336951237, 0.623251471203605, 1.23299690116447, -1.90252503712297, 
    -1.35720606056568, 8.07030264508413, 8.06895657403059, 8.07188495990973, 
    8.07156511986406, 8.0707792498515, 8.07413126898359, 8.06880946191224, 
    8.06797148880405, 8.06496363721434, 8.07013289455579, 8.07391287093536, 
    8.07358376989185, 8.07070251310967, 8.07103192180021, 8.07245964331964, 
    8.07244034544493, 8.07418273251513, 8.06811775036496, 8.0705566901228, 
    8.07071681967749, 8.06856533148604, 8.07134697455134, 8.06666030790906, 
    8.07020772302404, 8.06726582609184, 8.07372109797779, 8.06846181078564, 
    8.07259824748856, 8.07051451344483, 8.073172916069, 8.07359151970951, 
    8.06832275279002, 8.0744789611515, 8.07120733924244, 8.07155618881312, 
    8.07224977400496, 8.07448282679043, 8.06754100140664, 8.07697725917903, 
    8.07011751387304,
  0.0204912495149865, 4.92792788135823, 4.42892771485024, -3.51028368793088, 
    0.110792114307976, -0.503788987417965, 8.25406881108198, 
    -1.34417793845485, -2.79470932824448, -0.756018118105944, 
    8.80726715667119, 3.85061806713461, 1.67754461037642, 5.02909090726492, 
    1.36217748767801, -1.85834019268501, 1.76840303673449, 8.24484600503867, 
    -0.618407332735473, -4.81781850768985, -0.0144826471412252, 
    0.585082925398342, 2.1510458017186, 3.34557302677745, 5.64717135526349, 
    4.59706381568411, -2.87192791457713, 0.177768175998799, 1.91829401020921, 
    8.13802828397426, 6.34067258511198, -2.12741239410582, 
    -0.0709135699408986, 0.0350494091732371, 4.65437525028146, 
    8.48916173407804, 1.09637307793443, 1.21659517416449, -1.5454709452959, 
    -1.77407812359543, 8.03542041696532, 8.03407436953687, 8.03700275411904, 
    8.0366828456758, 8.03589704434403, 8.03924901332782, 8.03392726881541, 
    8.03308927731141, 8.03008139327377, 8.03525069933019, 8.03903064003953, 
    8.03870151748318, 8.03582028015038, 8.03614969095295, 8.03757736391871, 
    8.03755809792915, 8.0393004413899, 8.03323554525304, 8.03567438236178, 
    8.03583459353118, 8.03368307495765, 8.03646477561767, 8.03177814842985, 
    8.03532552057106, 8.03238359887089, 8.03883882600506, 8.03357956090628, 
    8.03771597426998, 8.03563231056605, 8.03829064202972, 8.03870928324275, 
    8.03344052476929, 8.03959675805874, 8.03632510799675, 8.03667397197315, 
    8.037367533488, 8.03960059382744, 8.03265881445794, 8.04209497637084, 
    8.03523525113418,
  -0.317212492661496, 4.97379236447749, 4.13635962633183, -3.7037320254914, 
    0.46254140300991, -0.184997435215918, 8.25326493359908, 
    -1.77567840947262, -2.97082078207585, -1.5317495430274, 8.48518272385518, 
    4.43050928780689, 1.18679106766224, 4.7794466885228, 1.89973040214864, 
    -1.81052900606636, 2.06278907478191, 8.00654868571635, 
    -0.0138104782106942, -5.27849936934571, -0.3156983342878, 
    0.825778079473971, 2.67114885115113, 3.26607945001906, 5.36826125939851, 
    4.90137446345955, -2.83497625790287, 0.153687628908648, 1.82546298520508, 
    8.04320458068236, 6.5476009887031, -1.98005212886339, 
    -0.0362400102718181, 0.115546547480747, 4.77017566353461, 
    8.42449874398598, 0.9427868315651, 1.14339208467743, -1.75525629177327, 
    -1.60846302249964, 8.06397430545092, 8.06262823591507, 8.06555663149028, 
    8.06523675046481, 8.06445091532022, 8.06780291626714, 8.06248111976788, 
    8.06164314035066, 8.05863527515481, 8.06380455500479, 8.06758451200612, 
    8.06725542370458, 8.06437416334577, 8.06470357190222, 8.06613127005658, 
    8.06611198350969, 8.0678543615251, 8.06178940687613, 8.06422830353564, 
    8.06438846641382, 8.06223698499115, 8.06501864248909, 8.06033198703543, 
    8.06387938302048, 8.06093748044152, 8.06739272777335, 8.06213343893068, 
    8.06626987749298, 8.06418616421115, 8.06684455788517, 8.06726316807608, 
    8.06199439617811, 8.06815061133675, 8.064878991286, 8.06522784571594, 
    8.06592142699551, 8.06815448368456, 8.06121266697818, 8.07064889170123, 
    8.06378915725283,
  -0.314359034880269, 4.99703006658665, 3.98685216753244, -3.72744357292166, 
    0.558939345345671, -0.182601283177884, 7.93722228421787, 
    -1.12283815671236, -3.22133333342956, -0.806402558256777, 
    8.83857334101238, 3.68937693690696, 1.57318758219653, 4.92145443163586, 
    1.5699797815566, -1.90072011535225, 1.90766581369581, 8.10022735762921, 
    0.288015641043651, -5.24674520004608, -0.266855695892704, 
    0.796421585641339, 2.38993686350013, 3.01497964498949, 5.28756218313998, 
    5.17209416242027, -2.65752123052182, -0.0642064195537139, 
    1.67985367193803, 7.89216462763377, 6.75095405777379, -1.88299122567471, 
    -0.205903829196005, 0.0775638762608419, 4.80330631182044, 
    8.35764130722934, 0.970940692001186, 1.18740292951605, -1.82217379904448, 
    -1.59580707840799, 8.02760110790151, 8.02625508359448, 8.02918345339096, 
    8.02886359655875, 8.02807774094011, 8.03142975208888, 8.02610794385596, 
    8.02526997627553, 8.02226210656555, 8.02743137672601, 8.03121136185529, 
    8.03088226536021, 8.02800100173359, 8.02833044361483, 8.02975815145291, 
    8.02973881964814, 8.03148124331796, 8.02541623414255, 8.02785519886498, 
    8.02801532380985, 8.0258638256226, 8.02864545825198, 8.02395876472847, 
    8.02750620468372, 8.0245643267701, 8.03101958196661, 8.02576027546353, 
    8.02989673840478, 8.02781301821873, 8.03047143532292, 8.03089003390867, 
    8.02562124204321, 8.03177747131575, 8.02850581414841, 8.02885468793778, 
    8.02954826899491, 8.03178131317734, 8.0248395041164, 8.0342757372519, 
    8.0274159980737,
  0.117519311651191, 5.46739030536232, 3.34809026894913, -3.72101431181503, 
    0.593190470361964, -0.0106573413657495, 7.5664883154404, 
    -0.800208012155097, -3.42160828179405, -0.544471121666457, 
    8.85272400087381, 3.55388092738235, 1.66835552623124, 4.96624101676011, 
    1.56416898239133, -1.8816198928808, 1.92208159468453, 8.00038616173523, 
    0.0757325820949601, -5.05870368197023, -0.0521556254093503, 
    0.523941847749867, 2.05671462441274, 3.28293306617463, 5.71520404959678, 
    4.5465824631255, -2.86568377906143, 0.200183609130645, 1.99225340835735, 
    8.17338643572683, 6.3584164500784, -1.99656853717079, -0.1027961459836, 
    -0.0194602942839972, 4.55433168975101, 8.54163979457054, 
    1.16066335809034, 1.25075879505238, -1.30513956545727, -1.73971193541909, 
    7.95918367103545, 7.95783760414266, 7.96076599155856, 7.96044613700808, 
    7.95966028400021, 7.96301228327824, 7.95769049669271, 7.9568525126037, 
    7.95384466553333, 7.95901392696922, 7.9627939097746, 7.96246480228944, 
    7.95958353960479, 7.95991293241274, 7.9613406532126, 7.96132136108732, 
    7.9630637497179, 7.95699878358154, 7.95943770781534, 7.95959783838415, 
    7.95744635293372, 7.96022799934616, 7.95554134415352, 7.95908875036341, 
    7.95614684751349, 7.96260212301442, 7.95734284239465, 7.96147925410342, 
    7.95939553922897, 7.9620539339094, 7.96247254083575, 7.95720377895939, 
    7.96335998469853, 7.96008836271643, 7.96043721561093, 7.9611307978873, 
    7.96336384691074, 7.95642203654687, 7.9658582785251, 7.95899852959397,
  -0.276440416809031, 5.37283211470841, 3.32109435950181, -3.86114642484759, 
    0.724475040860874, -0.0287271442330769, 7.69393242470942, 
    -0.729442309362226, -3.56699878084614, -0.588416339871392, 
    9.02452986806081, 3.35842501592024, 1.60792201177283, 4.96436232960491, 
    1.7388405796156, -1.89742403475109, 2.02773432757523, 7.98145948360863, 
    0.30889271189946, -5.17369923147168, -0.229193358958624, 
    0.58698268918155, 2.23682654392546, 3.06408841259125, 5.33702729205539, 
    5.0920723540179, -2.62915577974353, -0.0303953731153453, 
    1.76514278278224, 8.11056033696878, 6.22164020229642, -2.31497623452253, 
    -0.0219635463758729, 0.0614664387453267, 4.66419209312795, 
    8.45236110518982, 0.969404038738555, 1.17600559940111, -1.59172215559773, 
    -1.652597119768, 8.00738277639191, 8.00603672867529, 8.00896510508054, 
    8.00864522913353, 8.00785939542875, 8.0112113819052, 8.00588960376911, 
    8.00505162086688, 8.00204375664855, 8.00721305279792, 8.01099299504794, 
    8.01066389448806, 8.00778263831224, 8.00811205431282, 8.00953974857633, 
    8.00952047432461, 8.01126282626436, 8.00519790064347, 8.00763678512729, 
    8.00779695804257, 8.00564545608107, 8.00842712947837, 8.00374047127462, 
    8.0072878664228, 8.00434594467898, 8.01080120198173, 8.00554193083171, 
    8.00967835251826, 8.00759465964109, 8.01025302978231, 8.01067164434938, 
    8.00540288796691, 8.01155910668239, 8.00828746322321, 8.0086363405547, 
    8.00932990211268, 8.01156295088977, 8.00462114903276, 8.01405735977919, 
    8.00719763697448,
  -0.12986149978849, 5.25835687042205, 3.61251092582236, -3.81316439942048, 
    0.579302069401184, -0.183043707147095, 7.89968365596522, 
    -1.1848369128114, -3.54073052415024, -1.09894087768424, 8.66802830082722, 
    3.5727825986866, 1.25840179379614, 4.81843299469065, 2.70240068033118, 
    -1.77352215604435, 2.42714553405338, 7.74579833332005, 0.758103249909387, 
    -5.29193588944749, -0.153377055371735, 0.720388869312733, 
    2.18080120319355, 2.97510797339549, 5.36465045888181, 5.12905693343987, 
    -2.70698061522035, 0.00497131476533778, 1.88516700332878, 
    8.17833155718081, 6.32904132744633, -1.77764387645256, 
    -0.102127333566542, 0.0896917595409188, 4.72331231373081, 
    8.39870625540292, 1.03122987675872, 1.25666541551762, -1.56487301255743, 
    -1.68217851585244, 8.00741530401534, 8.0060692253455, 8.00899758785669, 
    8.00867773464134, 8.00789190994912, 8.01124392436385, 8.0059220863192, 
    8.00508413675201, 8.002076265909, 8.00724558230377, 8.01102551552927, 
    8.01069643539476, 8.00781516196893, 8.00814457366972, 8.0095722980159, 
    8.00955299960718, 8.01129534944308, 8.00523038727878, 8.0076693259108, 
    8.00782947167694, 8.00567797455919, 8.00845961002119, 8.00377297672134, 
    8.00732036584133, 8.00437846873255, 8.01083376277377, 8.00557443325641, 
    8.00971088695568, 8.00762716033118, 8.0102855403873, 8.01070416441206, 
    8.00543538345442, 8.01159164291014, 8.00832000677415, 8.00866885301168, 
    8.00936240635865, 8.01159548137271, 8.00465364914205, 8.01408991299112, 
    8.00723018592259,
  -0.139874137453125, 5.06768012294127, 3.98642904519815, -3.6637988603706, 
    0.465124673262024, -0.0973597399592421, 8.10466004064337, 
    -1.47889301655387, -2.943288884351, -0.985492244241175, 8.65659860348103, 
    3.91460840835776, 1.34623513939264, 4.79639635066083, 1.77194495009804, 
    -1.94183325839321, 1.90697107666205, 8.03136556143984, 0.422727490421621, 
    -5.00373816148072, -0.0180834356524149, 0.386195042802384, 
    1.74573820809617, 3.03142238599138, 5.6796698651692, 4.69169917554114, 
    -2.99135897847124, 0.196263526535561, 1.86068570261574, 7.98480666619069, 
    6.4175731439565, -2.04352110427575, -0.143421534203664, 
    0.0253022430945165, 4.62930540151735, 8.44405871810721, 
    0.994213163099299, 1.16113464844348, -1.55974766731165, 
    -1.61657630719968, 7.99949361091629, 7.99814755865982, 8.00107593428089, 
    8.00075607634159, 7.99997023660818, 8.00332223050347, 7.99800043863826, 
    7.9971624619185, 7.9941546085506, 7.99932388139336, 8.00310385230915, 
    8.00277475151378, 7.99989348660693, 8.00022289117271, 8.00165061057424, 
    8.0016313036325, 8.00337369823024, 7.99730872736595, 7.99974765495288, 
    7.9999077936817, 7.99775629845314, 8.00053793545643, 7.99585128569006, 
    7.9993986989615, 7.99645679426053, 8.002912074556, 7.99765278400758, 
    8.00178920272798, 7.99970549054309, 8.00236387584451, 8.00278249268421, 
    7.99751372687338, 8.00366994500814, 8.00039830862238, 8.00074717038143, 
    8.00144074830655, 8.00367378744328, 7.99673198092656, 8.00616822296946, 
    7.99930847707628,
  -0.262525520918977, 5.13359148852163, 3.78241097546787, -3.76902596065026, 
    0.621931928169215, -0.0219989189485225, 8.19881738600059, 
    -1.64821894891131, -3.16301254772614, -1.32255359063362, 
    8.62141709764742, 4.26670662308063, 1.35069678922176, 4.78220837628817, 
    1.55941552491272, -1.88987200016736, 1.86082621795107, 7.97663478736867, 
    0.290240019351574, -5.16355716592883, -0.106957004760248, 
    0.69901555636597, 2.15741582669857, 3.27323145673658, 5.80584345098857, 
    4.51179498477591, -3.00559405118549, 0.411426876579155, 2.28054261615895, 
    8.45961935509753, 6.10732834559132, -1.94234069393831, 0.145221483014571, 
    0.248241688964445, 4.86600114276714, 8.4329041761992, 0.80460601712714, 
    1.20178599029074, -1.56421233569485, -1.60210956416294, 8.00839826825927, 
    8.00705220350632, 8.00998058051552, 8.00966071819126, 8.00887488620766, 
    8.01222688635793, 8.00690508884949, 8.00606710769461, 8.00305924704091, 
    8.00822855013755, 8.01200847646248, 8.01167938758734, 8.0087981356615, 
    8.00912754639362, 8.01055525641482, 8.01053595792995, 8.01227831922102, 
    8.00621337721533, 8.00865227291124, 8.0088124356927, 8.00666095661982, 
    8.00944259275307, 8.00475595679702, 8.00830335169671, 8.00536144905837, 
    8.01181671527614, 8.00655742523597, 8.01069385001121, 8.00861015792448, 
    8.01126849166248, 8.0116871300951, 8.0064183616785, 8.01257461341454, 
    8.00930296502467, 8.00965182197099, 8.01034538878904, 8.01257843691073, 
    8.00563662630269, 8.01507286386549, 8.00821313730201,
  -0.518768345286787, 4.51239685524575, 4.27333625494237, -3.75673383270087, 
    0.914015163789295, 0.100089336583331, 7.75827894691075, 
    -1.24223688806902, -3.24490732744568, -1.14120284967014, 
    8.60469206355597, 3.83279169501874, 1.34714937774136, 4.90669421561479, 
    2.15746217664839, -1.8928714069162, 2.15672301512629, 7.96950998389347, 
    0.103710293363436, -5.11008239034809, -0.0343807464256609, 
    0.453121181048804, 2.09214286837678, 3.50037276416095, 5.92472046391201, 
    4.12508692889194, -3.05253553536386, 0.366342593604163, 2.06367460701728, 
    8.23734435930105, 6.46645933650907, -2.18391907238482, 
    0.0646766565813522, 0.248457225907412, 4.97377469379625, 
    8.31254671756302, 0.561297745405431, 0.999830070519789, -2.0685797772306, 
    -1.21041270502887, 8.03150179781895, 8.03015575450017, 8.03308413936285, 
    8.03276424381922, 8.03197842505561, 8.03533041591577, 8.03000865225814, 
    8.02917067056662, 8.02616277999127, 8.03133207474173, 8.03511201242609, 
    8.03478289442002, 8.03190165985302, 8.03223108296755, 8.03365877255573, 
    8.03363947936692, 8.03538184588343, 8.02931693073963, 8.03175576911166, 
    8.0319159826211, 8.02976447510715, 8.0325461500133, 8.02785951436768, 
    8.03140691492515, 8.02846497738709, 8.03492021666986, 8.02966094713014, 
    8.03379738094535, 8.03171369793308, 8.03437202256843, 8.03479066986187, 
    8.02952191401013, 8.03567813418865, 8.0324065017229, 8.0327553503427, 
    8.03344894126259, 8.03568197242455, 8.02874019014424, 8.03817637890723, 
    8.03131664939947,
  -0.524247091537664, 4.81042985711354, 4.06804698960163, -3.73892386867172, 
    0.657322944039983, 0.0829185093234054, 8.08270285514388, 
    -1.47214876998365, -3.15547407928472, -0.957973234992209, 
    8.74899110773033, 3.93427774740379, 1.40756822883404, 4.78063040122583, 
    1.67087417137619, -1.86348474999147, 1.92986133088177, 8.04771196462836, 
    0.259731718134866, -5.27920765345308, -0.274535477205888, 
    0.929250897409385, 2.42036715900143, 3.00155199753099, 5.30395026152006, 
    5.10898551975184, -2.69315788934381, 0.0368829519513042, 
    1.87809595364501, 8.14943258994377, 6.10707020967438, -2.05866492165148, 
    -0.0383035327879134, 0.131496777036977, 4.67387816745871, 
    8.39581740346652, 0.835081730962566, 0.910333088382922, -1.8459603681562, 
    -1.49926563994531, 7.99216069638106, 7.99081462203453, 7.99374300855119, 
    7.99342312325948, 7.99263730139026, 7.99598928957785, 7.99066750620387, 
    7.98982952286808, 7.98682166668538, 7.99199096684712, 7.99577095613208, 
    7.99544182970227, 7.9925605557661, 7.99288994647633, 7.99431765513644, 
    7.99429837990367, 7.99604074514278, 7.98997580240476, 7.99241472110015, 
    7.99257483699697, 7.99042337023847, 7.99320500570653, 7.98851837392195, 
    7.99206576051973, 7.98912385547071, 7.99557914645515, 7.99031984208715, 
    7.99445625499756, 7.99237255762054, 7.99503095324042, 7.99544954929001, 
    7.99018080044662, 7.9963370203659, 7.99306537154403, 7.99341423299669, 
    7.99410780012541, 7.99634086335412, 7.98939905234375, 7.99883529832211, 
    7.9919755489683,
  -0.226323034565638, 5.0976101033251, 3.74264678470129, -3.80124320782787, 
    0.691450053668973, -0.0231791575212523, 7.84645118821238, 
    -1.03576689100415, -3.48541811446948, -0.848713345419643, 
    8.91996299087429, 3.69443293573235, 1.48417803452158, 4.87525474338541, 
    1.66164977875425, -1.89473057017114, 1.92318346013574, 8.03583073788197, 
    0.206388058344528, -5.12385405399042, -0.11677363186559, 
    0.583701797856852, 2.09978112329911, 3.1447023114882, 5.58463341576214, 
    4.84964985763133, -2.81191625576819, 0.163817783267612, 1.91874465515027, 
    8.20178914839305, 5.89922720343896, -2.4884868226456, 0.191180297020258, 
    0.228478900269792, 4.72074386750723, 8.42611477448161, 0.867820972790725, 
    1.04326212266515, -1.54893915527809, -1.64931483896053, 8.00782376952714, 
    8.00647769059994, 8.00940609007054, 8.00908622063119, 8.00830038646785, 
    8.01165236997957, 8.00633058504877, 8.00549260580793, 8.0024847561502, 
    8.00765401387914, 8.01143402550807, 8.01110490122478, 8.00822363277132, 
    8.00855302872256, 8.00998075260065, 8.00996145004056, 8.01170385694865, 
    8.00563886861686, 8.00807781078869, 8.0082379249248, 8.00608645435083, 
    8.00886809053796, 8.00418142609625, 8.00772883661468, 8.00478695151917, 
    8.01124221926609, 8.00598293279347, 8.01011935152001, 8.00803563027864, 
    8.01069404545936, 8.01111263588265, 8.00584388302147, 8.01200007727996, 
    8.00872845741806, 8.00907730590392, 8.00977089174689, 8.01200394288698, 
    8.00506214409099, 8.0144983727128, 8.00763862753318,
  -0.299584307792025, 4.7658835773, 4.07448529476109, -3.69354501014783, 
    0.731993821913461, 0.159049140135372, 7.98486280647756, 
    -1.66270292890409, -3.06633925455477, -1.17511313238765, 
    8.48973498103957, 4.04216806729549, 1.31488651319543, 4.75493060541486, 
    2.01950852438473, -1.85851533623914, 2.07675981617454, 7.83744155600707, 
    0.62894522434175, -5.30416527742944, -0.130705484472634, 
    0.774188231234719, 2.18274145197048, 2.91652942289733, 5.2834665741847, 
    5.24104419360884, -2.59818669531973, -0.0699248761988281, 
    1.87028711943032, 8.36866531825977, 6.25105702112905, -2.11013303998433, 
    -0.0567528976182276, 0.161432958449411, 4.89530859272948, 
    8.42166300000378, 0.610990452098406, 1.18909680087774, -1.72839641184089, 
    -1.38660234962718, 7.96687979380535, 7.96553371778864, 7.96846211495534, 
    7.96814225944759, 7.967356405646, 7.97070839979865, 7.96538659893479, 
    7.96454862188107, 7.96154078042311, 7.96671003639674, 7.97049000646935, 
    7.97016090934005, 7.96727964758088, 7.96760904698698, 7.96903675792876, 
    7.96901746397679, 7.97075985519893, 7.9646949054728, 7.96713381793333, 
    7.96729393636433, 7.9651425002363, 7.96792412049282, 7.96323745686687, 
    7.96678486700542, 7.96384296740645, 7.9702982302108, 7.96503894401113, 
    7.9691753610839, 7.96709166403849, 7.96975004917274, 7.97016864693807, 
    7.96489990018165, 7.97105608835623, 7.96778446505078, 7.96813333303679, 
    7.96882692768892, 7.97105994602706, 7.96411814711092, 7.97355438203183, 
    7.96669464576078,
  -0.113945731981025, 5.43587732994441, 3.33117531094438, -3.81780654258476, 
    0.700605136059445, -0.0536140523688248, 7.76575233289434, 
    -1.09369986050594, -3.38349121041892, -1.01733098608725, 
    8.82132886856478, 3.86276294923876, 1.49533292982376, 4.94226820543944, 
    1.72454629561136, -1.88409613637066, 2.0017134701908, 8.02895379871278, 
    0.166178194653792, -5.11374270166583, -0.13126986785241, 
    0.645735506286842, 2.22632672477898, 3.31116430897289, 5.69577417443581, 
    4.50365018652065, -2.98007399626251, 0.369315547670019, 2.12162815977493, 
    8.22353660956718, 6.30146537432365, -1.92353816247988, 
    0.0033470270508455, 0.089547340715448, 4.69158650515017, 
    8.50017982085899, 1.01040746609865, 1.20642329469223, -1.47938940107115, 
    -1.6041310747777, 8.08551297125889, 8.08416690961867, 8.0870953080181, 
    8.08677544038378, 8.08598959009839, 8.08934157935975, 8.08401981061151, 
    8.08318183786841, 8.08017397070131, 8.08534321992756, 8.08912321426503, 
    8.0887940709429, 8.08591282021854, 8.08624222918952, 8.0876699560028, 
    8.08765064186004, 8.08939303964304, 8.08332810735847, 8.08576698612182, 
    8.08592712957162, 8.08377567563915, 8.08655729087391, 8.08187063819711, 
    8.08541805927601, 8.08247613915542, 8.08893140440042, 8.08367213772778, 
    8.08780856099977, 8.08572486657001, 8.08838322215175, 8.08880183856545, 
    8.08353311357765, 8.08968927367091, 8.08641766165213, 8.08676650376457, 
    8.08746012017125, 8.08969311101182, 8.08275134440386, 8.09218756434326, 
    8.08532783705433,
  -0.304686581743721, 5.09572631917949, 3.89180524490861, -3.74292568104153, 
    0.521012960571649, -0.0590072543646425, 8.14452799946953, 
    -1.36063445185199, -3.3270346377519, -0.945856332970652, 
    8.80041313134136, 3.81975658780775, 1.46558560321401, 4.85167783922558, 
    1.53850996122419, -2.05162262833551, 1.79982051386106, 7.97742584466426, 
    0.711923185851726, -5.22670146081735, -0.08878816940969, 
    0.451278572436922, 2.06240084173674, 3.05069378241207, 5.3132067225937, 
    4.81936647741242, -2.97307691772225, 0.170593476283579, 1.73798863941954, 
    7.91940186164511, 6.83136584001506, -1.51011645556042, 
    -0.106193674661637, 0.0865075334673231, 4.70457082578964, 
    8.38530287835568, 1.09682127669, 1.09124053017344, -1.74124087587041, 
    -1.5834623024186, 8.01807936325379, 8.01673331460977, 8.01966171025855, 
    8.01934182752001, 8.01855597683289, 8.0219079718343, 8.01658621142287, 
    8.01574822406507, 8.01274035630668, 8.01790962531373, 8.02168960083637, 
    8.02136048366171, 8.01847923510808, 8.01880864152949, 8.02023634567571, 
    8.02021706158303, 8.02195943955294, 8.0158944865203, 8.01833337451123, 
    8.01849354344846, 8.01634204058426, 8.01912370343061, 8.01443704978646, 
    8.0179844480531, 8.01504253840339, 8.02149779501299, 8.01623852535071, 
    8.02037495554641, 8.01829123457567, 8.02094963985784, 8.02136824542017, 
    8.01609948406845, 8.02225567745636, 8.01898405306764, 8.01933291706058, 
    8.02002650011052, 8.02225954037359, 8.015317730937, 8.02475396079352, 
    8.01789421744061,
  -0.173230665310157, 5.00314419543503, 3.9502198996633, -3.65032349302177, 
    0.573564137505189, -0.0793812476320124, 8.18629072165026, 
    -1.60072521404298, -2.96096175398407, -1.4212303582973, 8.55858647544619, 
    4.56054968380999, 1.13849378589207, 4.70472221145349, 1.18910338679619, 
    -1.82365217249095, 1.29774367644522, 8.45946343535243, 
    -0.685806504964801, -4.52482181001072, 0.405723865133667, 
    0.645020576748077, 1.72172493182298, 3.06257084653963, 5.65500752124025, 
    4.8633244561718, -2.7216686783332, -0.00487478829395407, 
    1.91236143233994, 8.17995563539584, 6.42313102150695, -1.77777165481853, 
    -0.175478686230646, 0.0946266202037002, 4.80149376781209, 
    8.41764776962952, 0.905075976205671, 1.24922507848941, -1.61512222166897, 
    -1.52730766806292, 7.92336688805632, 7.92202085401036, 7.92494924127607, 
    7.92462936309996, 7.92384350864419, 7.92719550110342, 7.92187374576224, 
    7.92103576056517, 7.91802789329381, 7.92319715520916, 7.92697712184849, 
    7.92664800914275, 7.92376676157872, 7.92409617103239, 7.92552387803148, 
    7.92550458445991, 7.92724695889491, 7.92118202736083, 7.92362090171462, 
    7.92378107696411, 7.92162957308675, 7.9244112248784, 7.91972458097954, 
    7.92327198192452, 7.92033006270417, 7.92678532629286, 7.92152606082778, 
    7.92566248068032, 7.92357878288599, 7.92623714909013, 7.92665577907829, 
    7.92138701825894, 7.92754321734178, 7.92427157960517, 7.92462045034877, 
    7.92531403000848, 7.92754704809312, 7.92060526203534, 7.93004148470833, 
    7.92318174987427,
  -0.40115777056715, 4.92052563413108, 3.87225369872778, -3.83580477853316, 
    0.841725113555308, 0.0674019767312087, 7.88556539897793, 
    -0.941035942622286, -3.40997106627307, -0.695695192510172, 
    9.02545700481161, 3.49253027413176, 1.56188160588596, 4.98344481443222, 
    1.77007624270776, -1.8625633175216, 2.0519896353915, 8.07039510444982, 
    -0.139993583052757, -5.13323131625126, -0.289671211074301, 
    0.712159542475445, 2.2036495549443, 2.90141376729569, 5.20633887922412, 
    5.36014982693967, -2.58257789067336, -0.10689931604196, 1.85127286854861, 
    8.47738313438564, 6.20591656087827, -1.98335862250933, 
    0.0809093686509532, 0.243268506423835, 4.96635325863434, 
    8.36531669216762, 0.638819492812426, 1.22676671874763, -1.82255398981458, 
    -1.41426404570477, 8.06846234170185, 8.06711628915093, 8.07004470604068, 
    8.06972480342422, 8.06893895001756, 8.07229094089575, 8.06696919470407, 
    8.06613120397202, 8.06312333108995, 8.06829258978862, 8.07207257597708, 
    8.07174344634829, 8.06886219335666, 8.0691915973078, 8.07061930370594, 
    8.07060002039775, 8.07234240468507, 8.06627747839485, 8.06871632417866, 
    8.06887650714802, 8.06672502587645, 8.0695066754376, 8.06482002607393, 
    8.06836743231951, 8.06542549066054, 8.0718807533012, 8.06662149956331, 
    8.07075792433245, 8.06867421751179, 8.07133259636741, 8.07175120496822, 
    8.06648247300766, 8.07263863105287, 8.06936702434204, 8.06971587652308, 
    8.07040948850625, 8.07264249401368, 8.06570070752615, 8.07513693919375, 
    8.06827719695996,
  -0.228493532511315, 4.01266826710034, 4.90070103787281, -3.42350001443195, 
    0.569169234125315, -0.23636465842612, 7.93171234936908, 
    -1.11379300006311, -3.24972949034449, -0.718952007038176, 
    8.78042222681452, 3.75706213423591, 1.65081940053054, 4.88567838171005, 
    1.42679232120105, -1.88735005160881, 1.84716047516235, 7.97798744964829, 
    0.205638730648277, -5.11515690617655, -0.0999123324620407, 
    0.61734485359874, 2.0070715963771, 3.23421587966523, 5.88122608658116, 
    4.56929822399671, -3.05688901051128, 0.224979426012832, 2.19232803904873, 
    8.01139660467329, 6.7239896531701, -1.06354423478938, -0.552630384544409, 
    0.167867212212942, 5.07090709328174, 8.290340094563, 0.381796170999979, 
    1.10261271535382, -2.11497564803304, -1.1378316898296, 7.98823551735857, 
    7.98688944912851, 7.9898178374436, 7.98949798195226, 7.98871213211933, 
    7.99206412451703, 7.98674233420945, 7.98590435359436, 7.98289651080578, 
    7.98806577161356, 7.99184575888971, 7.99151665363652, 7.98863538649759, 
    7.98896478319789, 7.99039250230641, 7.9903732077793, 7.99211559811532, 
    7.98605062448719, 7.98848956566684, 7.98864968067168, 7.98649820360497, 
    7.98927984174456, 7.98459318188966, 7.98814058577295, 7.98519869800208, 
    7.99165397209514, 7.98639468574395, 7.99053109914224, 7.9884473816722, 
    7.99110579368376, 7.99152439015991, 7.98625562927998, 7.99241183181391, 
    7.98914020093186, 7.98948906736043, 7.99018264016701, 7.99241568936382, 
    7.98547387732988, 7.99491011993895, 7.98805037529471,
  -0.347350816900127, 5.01593296587942, 3.80757071548226, -3.77757583547258, 
    0.749374612545308, 0.163793762919153, 8.027237597234, -1.52730496021347, 
    -3.13904417204666, -1.07976226073594, 8.77919135163033, 3.9809231864652, 
    1.46108817431654, 4.87446629490397, 1.63553067705725, -1.86674138672417, 
    1.94230198376834, 8.03684607779841, -0.038158653912507, -5.0913995204678, 
    -0.15892640702227, 0.629521948359716, 2.22623674074983, 3.19463308324997, 
    5.50040835762074, 4.87679033523887, -2.7695069413513, 0.0882558316037892, 
    1.90621231967459, 8.23731124056192, 6.17030572092168, -2.20736122309728, 
    -0.0201689204924612, 0.114272671510838, 4.66790638793541, 
    8.51051534479177, 0.750965136640775, 0.977914693239367, 
    -1.59973571382986, -1.48481311258288, 8.02392686230497, 8.02258079779885, 
    8.02550918787236, 8.02518927480246, 8.02440348565051, 8.0277554611353, 
    8.02243369602094, 8.02159570810946, 8.01858782515752, 8.02375714105605, 
    8.02753708337266, 8.02720796766652, 8.02432672951865, 8.02465615136156, 
    8.02608382480464, 8.02606454301798, 8.02780689388614, 8.02174196512274, 
    8.02418083548523, 8.02434101231636, 8.02218952674259, 8.02497119738521, 
    8.02028456967017, 8.02383194196727, 8.02089004743994, 8.02734528998544, 
    8.02208599904915, 8.02622242319896, 8.02413873729781, 8.02679709178197, 
    8.02721572064647, 8.02194696756458, 8.02810320639326, 8.02483154101686, 
    8.02518041701365, 8.02587396454196, 8.02810703296991, 8.02116522818688, 
    8.03060142216752, 8.0237416935017,
  -0.105412599749585, 5.28247748436679, 3.780864961269, -3.68229100522124, 
    0.42682794828759, 0.0147184876908682, 8.25172991542023, 
    -1.18102930481587, -3.37477737418256, -0.540214776166728, 
    8.84921541010917, 3.85869504943486, 1.55121541872458, 4.6456500392503, 
    1.08798022362243, -1.85780978847294, 1.54261115947275, 7.97331580068812, 
    0.271371237103, -5.24713797257452, 0.0284133930395608, 0.866975845802729, 
    2.00767181813475, 2.85522109647147, 5.44011062561969, 5.1051396948659, 
    -2.88025664893685, 0.174497106600831, 2.01994904867431, 8.28322074150722, 
    6.35976040920074, -1.6569236225783, -0.0346316128002389, 
    0.0871664644442532, 4.68061271624626, 8.50836423906896, 0.98653874205955, 
    1.23104063984162, -1.40444289654768, -1.66729810925408, 7.98221455819818, 
    7.9808684825776, 7.98379689319051, 7.98347701136312, 7.98269116346174, 
    7.98604316375959, 7.98072139007432, 7.97988342021203, 7.97687554193661, 
    7.98204479211434, 7.98582479724571, 7.98549565824022, 7.98261440722252, 
    7.98294381795856, 7.98437153293193, 7.98435223556912, 7.98609463027503, 
    7.98002967000896, 7.98246856216218, 7.98262871843162, 7.98047723461484, 
    7.98325888518668, 7.97857222790257, 7.98211963276152, 7.97917773135405, 
    7.98563297953098, 7.98037370113702, 7.98451014836057, 7.98242641694865, 
    7.98508483145329, 7.98550342642621, 7.98023468201667, 7.98639084534681, 
    7.98311924737477, 7.98346808342956, 7.98416169164944, 7.9863947264269, 
    7.97945292703947, 7.98888915080838, 7.98202940852029,
  -0.306482809433713, 4.94871332761196, 4.16861985500866, -3.65252358249977, 
    0.328187007639367, -0.349801049053413, 8.35859395538536, 
    -1.45875733855932, -3.20553457089926, -1.05380042611598, 
    8.72393895479729, 4.15833663716425, 1.52798395207237, 4.85128527836683, 
    1.30309887600045, -1.85507804707074, 1.71347283544741, 8.21000763284943, 
    -0.335320329089989, -4.83311085910646, -0.0620633067866272, 
    0.463704915638461, 2.02275957741672, 3.36088380191834, 5.7924508491995, 
    4.45498483413969, -2.88779704801822, 0.238173433621037, 2.09504962999805, 
    8.20260440395351, 6.40746293318597, -1.64614544976731, 
    -0.0669019653018174, 0.112452485595464, 4.78513217767121, 
    8.34808933120573, 0.98552021337187, 1.21447552255686, -1.79755397148235, 
    -1.64881752126976, 8.02952385738232, 8.02817777233927, 8.03110615371248, 
    8.030786323, 8.03000045552925, 8.03335247802775, 8.02803064959783, 
    8.02719267103568, 8.02418483699972, 8.02935411369169, 8.03313406247886, 
    8.03280498809332, 8.02992372285004, 8.03025311793485, 8.03168084837541, 
    8.03166155070173, 8.03340393156073, 8.02733894381565, 8.0297779004244, 
    8.02993800942638, 8.02778655071539, 8.03056816900372, 8.02588150983138, 
    8.0294289182045, 8.0264870251965, 8.03294231726361, 8.02768301386559, 
    8.03181944771473, 8.02973570638954, 8.03239411359034, 8.03281271169043, 
    8.02754394222129, 8.03370016151486, 8.03042854571256, 8.03077739820386, 
    8.03147097823223, 8.03370403190252, 8.02676218388561, 8.03619847034875, 
    8.0293387278312,
  -0.163283100324393, 4.78322549909868, 4.38842989243159, -3.56363476437656, 
    0.28589827162523, -0.207561969154715, 8.31929831071215, 
    -1.79003951477514, -3.00481367491899, -1.33987781013348, 
    8.51205619052662, 4.26526930494132, 1.04101653079694, 4.71325799396454, 
    2.44673198629728, -1.70503941429576, 2.28350781893976, 8.11184042471, 
    -0.379465415245936, -5.03557473484042, -0.260561033127615, 
    0.908132785178235, 2.18610625798584, 2.72255817779783, 5.03473973881781, 
    5.29366712296344, -2.83720341128218, 0.0614144128712611, 
    1.70137249731143, 8.08473913228813, 6.69997909489397, -1.47082365919798, 
    0.0852747165848475, 0.197528923980102, 4.78459790761426, 8.3182698412227, 
    1.02085139450423, 1.120318586731, -1.73551129536146, -1.66319718605868, 
    8.00287706406624, 8.00153097648397, 8.00445937684455, 8.00413954297176, 
    8.00335366977793, 8.00670566972681, 8.00138387770513, 8.00054589069197, 
    7.99753806094164, 8.00270730521189, 8.00648728921213, 8.00615818504279, 
    8.00327692205191, 8.00360630402944, 8.00503404021196, 8.00501474239139, 
    8.00675713877398, 8.00069217091875, 8.00313109833312, 8.00329120311518, 
    8.00113976213122, 8.00392137367569, 7.99923471272356, 8.00278212293363, 
    7.99984023268351, 8.00629551143791, 8.00103624161626, 8.00517264172678, 
    8.00308892310642, 8.00574731522911, 8.00616591430894, 8.00089716977661, 
    8.00705334960702, 8.00378174339924, 8.00413059413761, 8.00482418699776, 
    8.00705721537523, 8.00011539861511, 8.00955166181015, 8.00269192252411,
  -0.0825434983643389, 5.22147470659108, 3.76212697186415, -3.73661940218735, 
    0.591558967361238, -0.0171516767759521, 7.95779881782315, 
    -1.45819136085032, -3.2395402013826, -1.39760545648723, 8.73389973294814, 
    4.14313507015634, 1.20317313810874, 4.80220124919737, 1.75408668333671, 
    -1.88578716551245, 1.91479212443611, 8.01975763238024, 
    0.0619992066327909, -5.18437211851157, -0.144532303162586, 
    0.752053113267414, 2.21977124801726, 3.01117400363496, 5.351336115333, 
    5.15723025145894, -2.70292241039845, -0.0680873135395859, 
    1.74472147034637, 8.15181138622482, 6.62634416786979, -1.87882193785639, 
    -0.11499146429247, 0.0544989623889633, 4.68234564077275, 
    8.49757137023194, 0.996476683736807, 1.17102153682253, -1.47999805114547, 
    -1.65143638554943, 8.01542242370071, 8.01407640902919, 8.01700480255536, 
    8.01668492936499, 8.01589904682986, 8.01925104055345, 8.01392930498494, 
    8.01309131126572, 8.01008344645766, 8.01525268033441, 8.01903266331233, 
    8.01870353661589, 8.01582229818768, 8.01615169163719, 8.0175793910368, 
    8.01756011237849, 8.01930250690679, 8.0132375966441, 8.01567643567652, 
    8.0158366181673, 8.01368512606005, 8.01646678489163, 8.01178012461471, 
    8.01532753866472, 8.01238560294594, 8.01884083502237, 8.01358159573684, 
    8.01771801057733, 8.01563431898572, 8.01829272147501, 8.01871132868553, 
    8.01344256873424, 8.01959871811775, 8.01632711024588, 8.01667597810378, 
    8.01736960112829, 8.01960258951035, 8.01266080616901, 8.02209701415641, 
    8.01523726697171,
  -0.279204373550848, 5.45739864873271, 3.28325696275664, -3.84472266069634, 
    0.600198275887542, -0.067504904442334, 7.9307075051018, 
    -1.13022200969504, -3.48383334703006, -0.882751782498253, 
    8.8571937849543, 3.69359319436276, 1.42842524032945, 4.83937590325025, 
    1.88785367814308, -1.85664528609153, 2.05382021760152, 8.03493604906209, 
    0.301259482709976, -5.12252412841776, -0.222981534655274, 
    0.726825422567826, 2.07442590168288, 2.81481052440347, 5.22513905753157, 
    5.18075495519187, -2.73752740831676, 0.094146602438721, 1.87510823859013, 
    8.1668643974418, 6.42010571821944, -1.73090807521784, 
    -0.00985810547651953, 0.0938981877950675, 4.69502628592106, 
    8.37352720113264, 1.03677017723103, 1.22492690158734, -1.59253655664111, 
    -1.64831367098048, 7.97766161882506, 7.97631560454424, 7.97924396062344, 
    7.9789240648859, 7.97813826311855, 7.9814902411445, 7.97616848274155, 
    7.97533047696009, 7.97232259684892, 7.97749192859878, 7.98127181833487, 
    7.98094274035403, 7.97806150313845, 7.97839092970409, 7.97981858453639, 
    7.97979931416895, 7.9815416514909, 7.97547676776621, 7.9779155948066, 
    7.97807582002295, 7.97592429523859, 7.97870599835023, 7.97401936401471, 
    7.97756674930027, 7.97462482313774, 7.98108004385092, 7.97582077538544, 
    7.97995718190238, 7.97787355162642, 7.98053182755023, 7.98095050467852, 
    7.97568171716216, 7.98183800828301, 7.97856632085714, 7.97891520072118, 
    7.97960874079267, 7.98184181392211, 7.97490002924517, 7.98433618342897, 
    7.97747646732169,
  -0.0455608981647122, 5.13109707424141, 4.06071807578156, -3.74257936588567, 
    0.324414384898605, -0.22752116446022, 8.03234318191305, 
    -0.616672996939881, -3.72428367668268, -0.520227234097206, 
    8.78027301201107, 3.62036822261301, 1.39416669011879, 4.81639906596124, 
    2.07242584507777, -1.85626631569115, 2.19401534384603, 7.80934103860778, 
    0.6612087426094, -5.40582202500818, -0.256505725000193, 
    0.672208771349495, 2.674778091278, 3.4861447576816, 5.60501822001087, 
    4.83639782804135, -2.7208503740638, -0.00355373412047856, 
    1.83366946851941, 7.98591322417187, 6.54585064761594, -2.0677493034255, 
    -0.315428448532725, -0.0568990513363296, 4.5603122842627, 
    8.56352446004701, 1.04333638440616, 1.17654345385075, -1.398873783674, 
    -1.67319751974359, 8.07901509432209, 8.0776690623375, 8.08059745620858, 
    8.08027755215034, 8.07949171439101, 8.08284369677, 8.07752196206728, 
    8.07668396081779, 8.073676086867, 8.0788453684326, 8.08262530804923, 
    8.08229619984874, 8.07941496114127, 8.07974437542935, 8.08117205965925, 
    8.08115278568204, 8.0828951354017, 8.07683023510521, 8.07926906684092, 
    8.0794292770463, 8.07727776880543, 8.08005944485813, 8.07537281101228, 
    8.07892019523104, 8.07597825805805, 8.08243350675908, 8.07717425672825, 
    8.08131067294046, 8.07922699086301, 8.08188533072424, 8.08230397099474, 
    8.07703521692241, 8.08319142378952, 8.07991978040394, 8.08026865580903, 
    8.08096222788474, 8.08319525270502, 8.0762534707591, 8.08568966543311, 
    8.07882994341273,
  -0.110590706530969, 5.09628659278229, 3.83124022967111, -3.74781094625391, 
    0.619258974854021, -0.11765410462828, 8.03196541241656, 
    -1.54971375457014, -3.20637900593164, -1.41614931497804, 
    8.45071056143726, 4.54930040907244, 1.36963928381182, 4.77039995301078, 
    1.29916618319678, -1.95437258258884, 1.61059297681757, 8.20687916571864, 
    0.0149202028634183, -4.92208862840452, 0.0295367914548065, 
    0.448983695570298, 1.89938848047947, 3.13446625925814, 5.62213484715904, 
    4.81015087096294, -2.82184040725248, 0.07121802583826, 1.89243276943358, 
    8.0382850098146, 6.740406771654, -1.43697265484578, -0.228201915370721, 
    0.026899000446832, 4.65339183783144, 8.43024706942439, 1.04661033577912, 
    1.106739476791, -1.57803919400856, -1.50889452948294, 8.01148778760811, 
    8.01014174597292, 8.01307014589404, 8.01275026642317, 8.01196439029991, 
    8.01531640107932, 8.0099946288816, 8.00915664085512, 8.00614878546007, 
    8.01131804017365, 8.01509803162809, 8.01476892495089, 8.0118876585059, 
    8.01221705844644, 8.01364476385408, 8.0136254864972, 8.01536786867478, 
    8.00930292360386, 8.01174182020529, 8.01190196347817, 8.00975047964023, 
    8.01253211803434, 8.00784546586594, 8.0113928706037, 8.008450955199, 
    8.01490622545347, 8.00964694625182, 8.01378337391302, 8.01169966261427, 
    8.01435808225091, 8.01477667882858, 8.00950790947762, 8.01566409980726, 
    8.01239246410431, 8.0127413357271, 8.0134349272551, 8.01566795733674, 
    8.00872614413772, 8.01816240677364, 8.01130264852067,
  -0.537256197091065, 4.64564585233982, 4.26954025880738, -3.73349837047942, 
    0.620467621510845, -0.0824332048250613, 8.11380764310491, 
    -1.28250291282865, -3.28232368534472, -0.848898750283865, 
    8.8120109439833, 3.60149063963923, 1.4388370449108, 4.84236027054635, 
    1.95188714926856, -1.91237605265991, 2.08435793855097, 7.86260698386673, 
    0.646564755214852, -5.30194026446143, -0.182536512168, 0.697290600849214, 
    2.12711609802942, 2.93207802562815, 5.3484038565747, 5.15906653638385, 
    -2.62566455729648, 0.0272991275108649, 1.98272484083167, 
    8.28115168997947, 6.02269517065504, -2.07966565437261, -0.13162818576696, 
    0.0945302095556335, 4.79458880400817, 8.4127927046876, 0.657713026121688, 
    1.07896168668763, -1.97352197004489, -1.42236551110321, 7.98294558326362, 
    7.98159950713755, 7.98452792372909, 7.98420806390459, 7.98342218794943, 
    7.98677418864518, 7.98145241712395, 7.9806144301645, 7.97760658212024, 
    7.98277581094647, 7.98655581975426, 7.98622669276614, 7.98334544178605, 
    7.98367483882081, 7.98510255760049, 7.98508326157736, 7.98682567371404, 
    7.98076069839472, 7.98319960827185, 7.98335973195596, 7.98120827683735, 
    7.98398990694841, 7.97930323834344, 7.98285065326156, 7.979908758516, 
    7.98636401436958, 7.98110475223749, 7.98524117127287, 7.98315743789446, 
    7.98581586465371, 7.98623444653593, 7.98096570925892, 7.98712185660433, 
    7.9838502554555, 7.98419911438569, 7.98489272346629, 7.98712574295786, 
    7.98018392639904, 7.98962017732596, 7.98276042482702,
  -0.324209830308562, 5.29893235982138, 3.56485375499179, -3.82144192676757, 
    0.638266940318418, -0.114307182304105, 7.93150900464619, 
    -1.17192417181653, -3.33786261997368, -0.961945823672268, 
    8.82481768852127, 3.7457859238017, 1.51540013722363, 4.8819692592648, 
    1.54960974987328, -1.98715712415692, 1.83612971545542, 7.96099761827642, 
    0.745563554157423, -5.08206563688561, 0.013199661860015, 
    0.439376581782307, 1.64327927860511, 2.91873131061039, 5.79684223467347, 
    4.85289217939072, -2.9896828785113, 0.243280441163259, 2.12881442715077, 
    8.10264238759903, 6.55759787044778, -1.097988007609, -0.0837400461154813, 
    0.154399085280628, 4.75210605914477, 8.37047237756506, 1.09049283425813, 
    1.10556449558002, -1.70222873830406, -1.67028611821832, 8.02672420316288, 
    8.02537816018156, 8.02830652857939, 8.02798664235825, 8.0272008296428, 
    8.03055281415444, 8.02523103719566, 8.02439304562405, 8.02138518066587, 
    8.02655449737202, 8.03033444883051, 8.03000533881706, 8.02712407129747, 
    8.02745348847509, 8.02888118205474, 8.02886191433567, 8.03060426306148, 
    8.02453933305686, 8.02697822384767, 8.02713839142388, 8.02498687643591, 
    8.02776855898675, 8.02308190475666, 8.02662930783602, 8.02368737234463, 
    8.03014264864042, 8.02488336781179, 8.02901978504327, 8.02693609468487, 
    8.02959445932237, 8.03001307410705, 8.02474431911144, 8.03090056263414, 
    8.02762890474636, 8.0279777661494, 8.02867132438598, 8.03090439969854, 
    8.02396259874778, 8.03339880865806, 8.026539072337,
  -0.392499473229183, 5.0990764827088, 3.7720694924307, -3.78374303075138, 
    0.650395113433923, 0.0592489942430223, 8.23129800370934, 
    -1.71153781267895, -2.99045888847693, -1.20644721355831, 
    8.48853056952423, 4.24996523409565, 1.31139025966686, 4.79527492270146, 
    1.88620890934268, -1.87545998551872, 2.01090413999692, 8.14556847223393, 
    -0.0098633276177053, -4.90355028116298, -0.125149469424615, 
    0.340123620055077, 1.8471408695374, 3.33821951363625, 5.99423593390757, 
    4.41387387542748, -2.92861375150759, 0.280076371319442, 2.23697149454592, 
    8.30833431286358, 5.98224757853989, -1.85343409903402, 
    -0.0374838470069173, 0.144962178507639, 4.79533119393782, 
    8.38867909373199, 0.871548521324633, 1.19626544414008, -1.74128947085791, 
    -1.48979644240507, 8.0283539974413, 8.02700791325638, 8.02993631528084, 
    8.02961642788854, 8.0288305961077, 8.03218259893992, 8.02686079766677, 
    8.02602282343998, 8.02301495737478, 8.02818424413382, 8.03196425069274, 
    8.0316351323019, 8.0287538502456, 8.02908326262468, 8.03051096893227, 
    8.03049168840628, 8.03223406982247, 8.02616909505599, 8.02860802477236, 
    8.02876814601651, 8.02661667393632, 8.02939831565105, 8.0247116514068, 
    8.02825905685668, 8.02531716588032, 8.03177243902092, 8.02651313187588, 
    8.03064957630706, 8.0285658497039, 8.03122427553798, 8.03164285675212, 
    8.02637410176036, 8.03253031188588, 8.02925867775754, 8.02960752297614, 
    8.03030110210142, 8.03253418302501, 8.0255923585328, 8.03502861417188, 
    8.02816886370667,
  -0.406571004165805, 5.2263213739582, 3.59261158912344, -3.85072646376004, 
    0.740970672476169, 0.0122194957097221, 7.97956694175393, 
    -1.17680395142337, -3.33038578202609, -0.991475503398862, 
    8.97979971250576, 3.77395380312015, 1.51331248371588, 4.94511293007874, 
    1.30478299694581, -2.04459267198181, 1.62625405034601, 8.22108197820252, 
    0.47218751105086, -5.12163560634665, -0.0499594452105812, 
    0.712205542316377, 1.9717545195424, 2.77122923319316, 5.20495812281618, 
    5.2931442455368, -2.75912523937238, 0.0741544553406814, 1.75205225542562, 
    8.23547293677521, 6.43972895540232, -2.23495276129662, 0.1036726185819, 
    0.155497827486968, 4.78169193381622, 8.46006135576427, 0.798948637758606, 
    1.12800323323638, -1.6744859805859, -1.54853632189443, 8.06922667576122, 
    8.06788060559298, 8.07080901381003, 8.07048914261923, 8.06970329742369, 
    8.07305527754225, 8.06773352635354, 8.06689553824259, 8.06388767348669, 
    8.06905691358094, 8.07283689693617, 8.07250776670224, 8.06962652639311, 
    8.06995592916539, 8.07138364794331, 8.07136433702716, 8.07310673889628, 
    8.06704179832294, 8.06948066049591, 8.06964083249741, 8.06748936163197, 
    8.07027100304676, 8.06558435351936, 8.06913176367713, 8.06618985043712, 
    8.07264509390333, 8.06738584837319, 8.07152225741747, 8.06943856244958, 
    8.07209689668656, 8.07251553303787, 8.06724679834623, 8.07340296900008, 
    8.07013136827727, 8.07048020482664, 8.07117381096527, 8.07340682037463, 
    8.06646505294772, 8.07590124468317, 8.06904152433085,
  -0.606356044736804, 5.62647504569212, 2.99821453688666, -3.88763706191564, 
    0.733628162544898, 0.0242152465743451, 7.78291597018436, 
    -1.09810538716542, -3.41886684848707, -1.10708959953561, 
    8.83329629621015, 3.86342177927008, 1.55998237969649, 4.93907068151451, 
    1.23892839741974, -1.98515175566223, 1.67867281278768, 8.05320364942544, 
    0.381539133915975, -5.08597385857931, -0.0769596594931248, 
    0.474247206909897, 1.96104615991122, 3.13054981450627, 5.61836575358983, 
    4.67228088011472, -2.91920400014257, 0.27320377956501, 2.0090448434243, 
    8.09378636927625, 6.42539550420196, -1.6966465917576, 
    -0.0332049272290863, 0.0515550439733318, 4.63543582654365, 
    8.42915637014355, 1.09578679519818, 1.10984746349096, -1.73494254722875, 
    -1.49468574829189, 8.01730255787155, 8.01595651922586, 8.01888491223291, 
    8.01856502936031, 8.01777918300599, 8.02113117110105, 8.0158094239239, 
    8.01497143203498, 8.01196356354753, 8.01713282410434, 8.02091279593526, 
    8.02058366863244, 8.01770242414711, 8.01803182784637, 8.01945953567184, 
    8.01944024134609, 8.02118262259758, 8.01511770770499, 8.01755655798467, 
    8.01771673176534, 8.01556524921604, 8.01834689763547, 8.01366025687407, 
    8.017207661205, 8.01426572736656, 8.02072098765729, 8.01546173651436, 
    8.01959813724257, 8.01751445485402, 8.02017280764355, 8.02059143843127, 
    8.01532269271432, 8.02147887696076, 8.01820724747629, 8.01855611020167, 
    8.01924970742507, 8.02148271088946, 8.01454093499045, 8.02397714785256, 
    8.01711740773384,
  -0.290993581616183, 5.43863088372574, 3.2201779501282, -3.89281620189012, 
    0.726005525271891, 0.091650179639097, 7.73304722494163, 
    -0.675354867045794, -3.61771695357099, -0.512956606788042, 
    9.12680210781268, 3.51660626733362, 1.56821719111828, 4.9536783407016, 
    1.53715224160314, -1.82767738550953, 1.81584491080864, 8.28424885295201, 
    -0.398137328193538, -4.64856379488369, 0.0968458157734258, 
    0.444371424081891, 1.8283152339271, 3.29569738586288, 5.88428709615821, 
    4.37378593866186, -2.99618612999148, 0.241781517731152, 2.00758584551547, 
    8.20088568471901, 6.19251332623675, -2.09202053454323, 0.014317564337725, 
    0.130363065016649, 4.75386017196051, 8.39632604575926, 0.839222284351371, 
    1.25800132626391, -1.54834469152517, -1.60694817091808, 7.98863236093839, 
    7.98728629630161, 7.99021469920123, 7.9898948318532, 7.9891089736298, 
    7.99246096758681, 7.98713919775663, 7.98630121028669, 7.98329335435339, 
    7.98846261336477, 7.99224258530439, 7.99191346531101, 7.98903221877883, 
    7.98936162305795, 7.99078932864281, 7.99077004397935, 7.9925124244948, 
    7.98644748725843, 7.98888636780341, 7.98904651970801, 7.98689505395262, 
    7.98967669764544, 7.98499004184976, 7.98853744795931, 7.98559553645628, 
    7.99205078713132, 7.98679152299514, 7.99092794260387, 7.98884424058022, 
    7.9915026179166, 7.99192122295172, 7.98665248250128, 7.99280866315089, 
    7.98953704245597, 7.9898859011794, 7.99057949820029, 7.99281252321196, 
    7.98587072173291, 7.99530694872021, 7.98844721061204,
  -0.218810686770724, 5.06560353701816, 3.81042753361896, -3.77583788160221, 
    0.651783179408966, -0.118282933925343, 7.87325511943025, 
    -1.14343804018652, -3.32915460924096, -1.00694639236793, 
    8.84205353871546, 3.77985833975348, 1.38384921202435, 4.87834896567458, 
    1.89485672573845, -1.84811070388618, 2.05348392510215, 8.00809255204753, 
    -0.0535040176105584, -5.10097986729092, -0.177806402214942, 
    0.719986945759867, 2.15932888512659, 3.01470944220025, 5.40415058494694, 
    5.07241314699335, -2.72027774757266, 0.120702397005042, 2.05190864258728, 
    8.49225047669785, 6.28907741530787, -1.76892383612435, 0.128462619933979, 
    0.259318375214848, 4.92802926590092, 8.32785876372537, 0.777604868443965, 
    1.25295717137979, -1.67002867356168, -1.61560909004678, 7.98198321615522, 
    7.98063714515113, 7.98356555275457, 7.98324570230026, 7.98245984181191, 
    7.98581182211928, 7.98049005912308, 7.97965207884077, 7.97664422384279, 
    7.98181345617119, 7.98559345388438, 7.98526432399573, 7.98238307043508, 
    7.98271247337728, 7.98414021957949, 7.98412088915817, 7.98586332172298, 
    7.9797983289422, 7.98223723947102, 7.98239738235628, 7.98024591088148, 
    7.98302753483201, 7.97834086308615, 7.98188829096405, 7.97894638338533, 
    7.98540165542589, 7.98014240927929, 7.98427882330435, 7.9821950755891, 
    7.98485347783419, 7.98527207506642, 7.98000335337626, 7.98615948628177, 
    7.98288791310835, 7.9832367616348, 7.98393037466167, 7.98616336897862, 
    7.97922157172935, 7.98865780394908, 7.98179807424418,
  -0.322724286568128, 4.41740046156626, 4.82312184311829, -3.51674967837315, 
    0.306286948131109, -0.0522064746706552, 8.27551388227072, 
    -1.03318499162512, -3.48587932164866, -0.485274713348005, 
    8.86917390102343, 3.50841564324972, 1.52237111467643, 4.84053463001432, 
    1.76490354208103, -1.88205909651565, 2.02542755657853, 7.84653674472948, 
    0.621016084369699, -5.31178444740277, -0.163026788670183, 
    0.785297472369457, 2.34166613565224, 3.19624783241421, 5.56799056947405, 
    4.85782998124932, -2.77265744082977, 0.212686071160406, 2.18215938954828, 
    8.43568535954961, 6.27994890714895, -1.86828311571117, 
    -0.0914668756645965, 0.145794342143356, 4.88680121113695, 
    8.41775513635155, 0.612315789190401, 1.11260883708846, -1.86622438981741, 
    -1.33339027283214, 8.02739414416546, 8.02604809060182, 8.02897646755529, 
    8.02865658019538, 8.02787077484908, 8.03122274893747, 8.02590097389571, 
    8.02506299941621, 8.02205512303024, 8.02722443552378, 8.03100438403216, 
    8.03067525625705, 8.02779400303166, 8.02812342101152, 8.02955112289544, 
    8.02953182961647, 8.03127418817467, 8.02520927242348, 8.02764814474236, 
    8.0278083124659, 8.02565683241676, 8.02843847596914, 8.02375184094492, 
    8.02729923948168, 8.02435731979984, 8.03081258353943, 8.02555329752259, 
    8.0296897186895, 8.02760604555209, 8.03026437849087, 8.0306830064838, 
    8.02541426776777, 8.03157049413957, 8.0282988381347, 8.02864770115749, 
    8.029341273335, 8.03157430599683, 8.02463252530432, 8.03406873197025, 
    8.02720900830282,
  -0.305939533678084, 5.4418487892173, 3.22072677107858, -3.88573227306023, 
    0.741053549048193, 0.0944831146734445, 7.78973000286919, 
    -1.02508980194506, -3.62045736242677, -0.925394192907191, 8.908277916053, 
    3.56779428547674, 1.42561171784738, 4.88647066339301, 2.02471053407798, 
    -1.84678982780414, 2.13554683896162, 7.85741440235512, 0.422852582174117, 
    -5.26446327557875, -0.135001318947251, 0.779230492236235, 
    2.23366421395687, 2.99600598829399, 5.35094147585919, 4.95903412794035, 
    -2.93934202569759, 0.140887875492851, 1.79822850229907, 8.10929311396314, 
    6.56777908921737, -1.7323762466513, 0.0322114319428122, 
    0.176334885282822, 4.79089118106901, 8.37801128325349, 0.982863133123653, 
    1.19822160892355, -1.58731664062973, -1.6023199199457, 7.9875859683307, 
    7.98623992075608, 7.98916831045265, 7.98884842508051, 7.98806258763056, 
    7.99141456746643, 7.98609281119395, 7.98525482017367, 7.98224695822521, 
    7.98741622937332, 7.99119620030921, 7.99086708303036, 7.98798582983639, 
    7.98831523215649, 7.9897429227602, 7.98972364983505, 7.99146601702291, 
    7.98540110458539, 7.98783997127427, 7.98800013288208, 7.98584865116455, 
    7.98863031798416, 7.98394366601499, 7.98749105784182, 7.98454914057939, 
    7.99100438861699, 7.98574512539293, 7.98988152976958, 7.98779785227942, 
    7.99045622510152, 7.99087483863788, 7.98560608762467, 7.99176228271929, 
    7.98849064452103, 7.98883952068752, 7.98953309645268, 7.99176613097516, 
    7.9848243465878, 7.9942605427769, 7.98740080974075,
  -0.156921190290516, 4.9591290879662, 4.03135421000723, -3.75826202539549, 
    0.539156749778779, -0.151327454270928, 7.97416246653399, 
    -0.724916115756769, -3.59279472081216, -0.460689560376137, 
    8.96119342913155, 3.48965682580436, 1.50159088858115, 4.86540649682772, 
    1.79589459797696, -1.88608551119559, 1.98852028154303, 8.07362207050939, 
    0.0238090425239712, -5.03775813622008, -0.116231433965957, 
    0.477779511870783, 1.90786558074652, 3.03903767696992, 5.56134712394379, 
    4.93349287564284, -2.79293084813273, 0.110087429040359, 1.96616234452116, 
    8.33788403015794, 6.1649999980041, -2.06495274048926, 0.0542866330433486, 
    0.182856458551713, 4.86292267633949, 8.36822412358668, 0.841350548864406, 
    1.28535679915199, -1.64690912998263, -1.61803016202906, 8.00949634102645, 
    8.00815031405891, 8.01107870366186, 8.0107588263871, 8.00997297944187, 
    8.01332495590299, 8.00800322744853, 8.00716523328301, 8.00415735634677, 
    8.00932661481507, 8.01310654631992, 8.01277741574352, 8.00989620483992, 
    8.01022561121524, 8.01165329821088, 8.0116340050566, 8.01337638124143, 
    8.00731151194409, 8.00975030280635, 8.00991051612806, 8.00775904332965, 
    8.01054069997488, 8.00585406871434, 8.00940147235186, 8.00645952421944, 
    8.01291474611033, 8.00765551519382, 8.01179191236678, 8.00970826746163, 
    8.0123665553814, 8.01278521384624, 8.00751648131894, 8.01367265490405, 
    8.01040103162497, 8.01074989569065, 8.01144351202456, 8.01367648107086, 
    8.00673472972374, 8.01617089250929, 8.00931117137544,
  -0.636426774999669, 5.20604150871862, 3.39306074283717, -3.88899150454619, 
    0.858488546079597, 0.353036418520624, 8.01725224562311, 
    -1.30013691939824, -3.28770063435578, -0.628806298949203, 
    8.91593247691954, 3.4737045216091, 1.67911324895635, 4.96812058489155, 
    1.68540725737112, -1.86745279040382, 2.023737605285, 8.01927083955387, 
    0.362727961240916, -5.26284683925186, -0.256767285237787, 
    0.727578176560294, 2.5585650520198, 3.52586381734861, 5.73178267946263, 
    4.49694426102755, -2.83096575864115, -0.00494509051688862, 
    1.73278079079162, 7.5492464965112, 7.1134437522577, -1.14619705801904, 
    -0.540114245441576, -0.0346894798765593, 4.55051401144539, 
    8.39295360913508, 1.0418857272724, 0.807769817672887, -1.878423671483, 
    -1.29833489352635, 8.00088705065703, 7.99954097346399, 8.00246939276636, 
    8.00214951297082, 8.00136366151519, 8.00471565229355, 7.99939388911114, 
    7.99855590550956, 7.9955480389096, 8.0007172831151, 8.00449727104936, 
    8.00416813943424, 8.00128689814743, 8.00161629593959, 8.00304400782483, 
    8.00302471085572, 8.00476711357879, 7.99870216965446, 8.0011410284748, 
    8.00130119334625, 7.99914974346008, 8.00193137784696, 7.9972447246564, 
    8.00079213372301, 7.997850223362, 8.00430545853359, 7.9990461996675, 
    8.00318262378657, 8.00109891607409, 8.00375729541514, 8.00417590242598, 
    7.99890716602565, 8.00506332326996, 8.00179173127553, 8.00214057164045, 
    8.00283419355932, 8.00506720170521, 7.99812541109618, 8.00756162781606, 
    8.00070188844109 ;

 state_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1 ;

 state_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 time = 41.625 ;

 advance_to_time = 41.625 ;
}
