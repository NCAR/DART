netcdf filter_input {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 40 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;

	double state(time, member, location) ;
		state:long_name = "the ensemble of model states" ;

	double state_priorinf_mean(time, location) ;
		state_priorinf_mean:long_name = "prior inflation value" ;

	double state_priorinf_sd(time, location) ;
		state_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double state_postinf_mean(time, location) ;
		state_postinf_mean:long_name = "posterior inflation value" ;

	double state_postinf_sd(time, location) ;
		state_postinf_sd:long_name = "posterior inflation standard deviation" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "days" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id: $" ;
		:model = "Lorenz_96" ;
		:model_forcing = 8. ;
		:model_deltat = 0.05 ;
		:history = "identical (within 64bit precision) to ASCII filter_ics r1350 (circa June 2005)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 location = 0, 0.025, 0.05, 0.075, 0.1, 0.125, 0.15, 0.175, 0.2, 0.225, 0.25, 
    0.275, 0.3, 0.325, 0.35, 0.375, 0.4, 0.425, 0.45, 0.475, 0.5, 0.525, 
    0.55, 0.575, 0.6, 0.625, 0.65, 0.675, 0.7, 0.725, 0.75, 0.775, 0.8, 
    0.825, 0.85, 0.875, 0.9, 0.925, 0.95, 0.975 ;

 state =
  -2.072284116226430, 2.667234685046764, 5.544948506330924, 4.310057631263879,
    -1.669912120996396, 1.876109568728516, 6.097723157457765, 4.799036507527475,
    -4.988434568614633, 4.888450137598835, 5.305675918629604, 3.293790529508235,
    6.349049865798637, 4.014261196679387, 1.320815660634750, 3.965189184473605,
    2.678136186383346, -2.045969003028782, 2.213639991606812, 3.415866822965563,
    7.491227111954361, -2.536805899681665, -1.231290322654628, 1.581869564035022,
    3.255572179144334, 4.067728046168671, 5.763380760632609, -3.320369736559728,
    -0.4517825866222965, -1.764376279365341, 8.662830548905710, 1.644165971778301,
    1.553529010785091, 1.899340123523308, 3.579790688167297, 7.879578534281588,
    0.5974337791566716, 2.285632865564447, 5.664239076200905, 6.689938799827169,
  -3.202906134396487, 2.715681557300329, 5.108376283089062, 6.120608202038975,
    -0.6272239209739398, 1.245856523078123, 5.317388140041573, 6.401577193637829,
    -3.579996900491562, 5.866294219712250, 5.246267828512429, 2.022044006745020,
    5.848167914810999, 4.920581093177566, 1.019630791634363, 3.757669157386637,
    3.541050578368573, -1.964965359272030, 2.396254345729744, 3.723997890351967,
    7.433151081993870, -2.718570414603811, -1.223368863016383, 1.741714563075974,
    3.192490201334766, 3.778152136820833, 6.033810479676742, -3.294282828968004,
    -0.6111941274887129, -2.246927361835390, 8.606220419657969,
    1.725800163564966, 1.081262513612530, 1.650329356397879, 3.591284709413881,
    7.821704768816453, 1.027829743208568, 2.865344518372303, 6.401803040988903,
    5.233199003327673,
  -3.233288888140787, 2.791047456869411, 5.443532527304444, 5.271340589601074,
    -1.405216415938772, 1.865789062676320, 5.762713557048915, 6.180405666138984,
    -4.097543907249058, 5.423289545303277, 5.434883543884185, 3.005727493198202,
    6.145393134062668, 4.064569804715867, 1.341113924400163, 3.960643467935648,
    2.932665169142973, -2.104913189023151, 2.287547409452981, 3.578121373316026,
    7.512267541136903, -2.574491867576626, -1.366896665783236, 1.764350341552444,
    3.219368317877549, 3.762638146162343, 6.034752102196681, -3.336595117188780,
    -0.5646284297952464, -2.279574592228803, 8.536819705885497, 1.669626532010157,
    1.024001937708187, 1.671573610782606, 3.701025508503733, 7.828641074190320,
    0.8559438345358253, 2.727434162133096, 6.413964978404168, 5.530961064974001,
  -3.380206933377884, 2.905616122235494, 5.796544048481724, 4.762968769969448,
    -1.572686591853639, 1.992704930576504, 5.995706965663434, 5.629340431894160,
    -4.561161315439922, 5.226261209797866, 5.460717559795719, 3.069425527232305,
    6.173554911447423, 4.123680428751393, 1.145215572910912, 3.876153624231368,
    3.103547215145973, -2.085313305778273, 2.198468609227772, 3.233270352766603,
    7.826651493076933, -2.364471062614204, -1.236187695043357, 1.647284819778698,
    2.970635730634302, 3.718377516689948, 6.102637834877616, -3.253961411547286,
    -0.5740797521566847, -2.209320215434456, 8.657683346820132,
    1.673066851187036, 0.9653828495097909, 1.556198226880673, 3.517216765928562,
    7.959247064667264, 1.150916317449992, 2.797052145884083, 6.618709247272493,
    5.043448562643719,
  -3.407629759706746, 2.933433929830310, 5.866755154866184, 4.694034214784155,
    -1.501568595569831, 1.958730160918034, 5.993571164774017, 5.151337819723222,
    -4.944286584326520, 4.994702956954078, 5.236249746761420, 3.113257300241284,
    6.312305199725202, 4.360060672821684, 1.250993119716547, 3.873765648616770,
    2.802528892415240, -2.101359010997210, 2.087365453862844, 3.154883038801723,
    7.962039000133199, -2.335450842457444, -1.138455991039180, 1.604428995832406,
    2.840931890760030, 3.664057544364724, 6.169114960043840, -3.206745584619120,
    -0.5159824231897091, -2.139408571663462, 8.686732444575666,
    1.723929032670534, 0.9767155001336526, 1.545949842323754, 3.453550414329027,
    8.014161426610357, 1.263562428978997, 2.771743857242854, 6.592628223389382,
    4.895994327088172,
  -3.242250962223488, 2.963074836651538, 5.735156062293944, 4.956481603798761,
    -1.424562843101034, 1.912606251664502, 5.901836045695529, 5.717399776854215,
    -4.710704664707484, 5.124356898835035, 5.506509036254787, 3.524644752456478,
    5.796538782325586, 2.984026795105250, 1.615839609253615, 4.014968612172839,
    3.259495544690143, -2.135418016689775, 2.001809645421830, 2.202060531680972,
    8.358668976227230, -1.336194540907803, -1.603381151882028, 1.961111193267988,
    3.169038178219075, 3.711615245424609, 6.211766948247375, -2.903313512266379,
    -0.2636723127436703, -1.255774988255093, 8.934925759734595, 1.633322772458381,
    1.362774819919612, 1.625821482014907, 3.219348129773149, 8.154478543873864,
    1.519596200812855, 2.599593136279430, 6.377654226982051, 5.366944658663931,
  -3.362550518681563, 2.907490527111332, 5.754364141175526, 4.807819205952152,
    -1.524056795245456, 1.987058463913923, 5.929420671752847, 5.670521524704461,
    -4.598425379017116, 5.189115970890054, 5.389638923913724, 3.085457060774673,
    6.182833982228911, 4.135858704147793, 1.121602960366592, 3.854968884980818,
    3.133874700525292, -2.066803878799485, 2.186409174498391, 3.124928762295082,
    7.862155379129307, -2.284354407552081, -1.249830410826104, 1.639642006679358,
    3.009739683109256, 3.784326284304012, 6.048564248069831, -3.257796017393361,
    -0.5372025103585109, -2.127954981734660, 8.713072883418535,
    1.627380651190578, 0.9453065559702664, 1.512906047829786, 3.443017925703078,
    7.967544104359317, 1.196063917869892, 2.814721319026404, 6.617711030292702,
    5.074171269337790,
  -3.294432115187644, 2.900818063554855, 5.671131525016277, 4.951869690302068,
    -1.521433928720328, 2.015400529692046, 5.999377166464523, 5.754511364452459,
    -4.250621279822100, 5.329718248513848, 5.635389989069359, 3.176689370084834,
    6.258560495972246, 4.316308337047451, 1.427463883454208, 3.900545151153008,
    2.506359015444425, -2.087468822618553, 1.982345742572358, 2.761460437266656,
    8.240171951600194, -2.039686303815361, -1.256206235532622, 1.711962537807816,
    2.938331749285644, 3.664040136850155, 6.177828482432234, -3.210410780259355,
    -0.6969942863679864, -2.256506320598111, 8.690814238420312,
    1.728772806801648, 1.108516822691623, 1.591829741951198, 3.484564977388727,
    7.887018825911350, 1.042085436028796, 2.768842579606509, 6.522307663121132,
    5.401230223832295,
  -3.469278631236071, 2.901890487693050, 5.570830379846906, 5.243372653072932,
    -1.167647118683344, 1.998459064929182, 5.862167678346749, 5.379212628999523,
    -4.803595272743691, 5.028353205580556, 5.404979899539868, 3.282237164426145,
    6.156517113129256, 3.829592217096554, 1.172766194102839, 3.882838637498282,
    3.223565615812178, -2.069594705868352, 2.160084183923471, 3.013183760043594,
    7.992015436745972, -2.168551775450724, -1.280567409665402, 1.721044157723455,
    2.996964488359199, 3.691880643221109, 6.132936771152680, -3.279198906460006,
    -0.5726429060047649, -2.228513566831877, 8.594570094660604, 1.758190723378030,
    1.096836293939859, 1.683480334481025, 3.674994312573483, 7.886592758448806,
    1.041958043202223, 2.809455140061428, 6.528615282141470, 4.834841980876813,
  -3.292301545328965, 2.965828151212683, 5.788344034308993, 4.869366231928398,
    -1.518652917279586, 1.885798171059188, 5.661007276886391, 6.309846061099589,
    -4.408874966864532, 5.179287402261099, 5.266935171059665, 3.216641304719170,
    6.099468101327123, 3.796293266161881, 1.135276712413784, 3.834357201868248,
    3.425784181446673, -2.114956063702472, 1.963212745571410, 2.661413710469108,
    8.402772169586573, -1.966250382809288, -0.8584614993121848,
    1.336424168821090, 2.332698275182698, 3.577264712695379, 6.266741809409380,
    -3.187908629758062, -0.2662083782113466, -1.584478708319061,
    8.487668144400795, 1.061265634828200, 0.8786507813482253, 1.673898765480351,
    3.882034754689747, 7.913696118795533, 0.8743563487025602, 2.642693771002228,
    6.452778989667022, 5.067159838828500,
  -3.131521665987826, 2.810929514637102, 5.473704591732365, 5.005860296467167,
    -1.520284429856362, 2.053959636186800, 5.854399607406782, 5.944804671598308,
    -4.321487887218949, 5.318028326371111, 5.188397052769758, 2.993001390004456,
    6.423473028579533, 4.857285017659472, 1.360719558438343, 3.725473527072056,
    2.122417993313940, -1.982210878403592, 1.982906428057667, 3.251425903547606,
    7.746590112937211, -2.470882577545793, -1.304372620932889, 1.683118926254431,
    3.071421656228133, 3.771927732178853, 6.135008715355539, -3.135117173751596,
    -0.6706897572540047, -1.916912940382090, 8.833271099521937,
    1.306474700199141, 1.047435745504077, 1.431426827655883, 3.171662889034394,
    7.985231731236074, 1.310136806078764, 2.632203335960277, 6.305108227159463,
    5.738298662267306,
  -3.090360605876935, 2.816398127961831, 5.342119240786285, 5.230074806145530,
    -1.215088731548626, 1.917815397371886, 5.762254538326108, 5.488829306692382,
    -4.908259737294575, 4.944970792786369, 4.866783676135982, 3.109029143631202,
    6.305561487670104, 4.200276191781060, 1.316676725476829, 3.866187116906347,
    2.907277141515618, -2.053437869037750, 2.006253123947553, 2.476595601574689,
    8.250432737800883, -1.755759431619256, -1.405818627989155, 1.807766363474797,
    3.105678640629238, 3.731821116456178, 6.071569463251309, -3.329647755145270,
    -0.5870743864176731, -2.352828452107243, 8.606144085239512, 1.745080051267500,
    0.9588852789408137, 1.562959656951018, 3.530027203180039, 7.816389267284324,
    0.8270604107103331, 2.733780265161935, 6.314456605151813, 5.813405496694255,
  -3.255438931889410, 2.874026591884559, 5.607949407292672, 4.947424226881743,
    -1.470559728530715, 2.006979814777722, 5.917301735320533, 5.678064496019751,
    -4.634524088589051, 5.169269416115695, 5.301418169628593, 3.129417629583326,
    6.239169318612233, 4.156938191770986, 1.220061519599440, 3.891634355740891,
    2.948702938576102, -2.065833363785824, 2.219763680080484, 3.230582878634644,
    7.789911870226623, -2.328416136530722, -1.358510049884152, 1.789819881985681,
    3.225853236466314, 3.788601474935912, 6.035080364570865, -3.312914433355886,
    -0.5760426032409967, -2.240456823633295, 8.618080323437216,
    1.745338699233793, 1.067137650957099, 1.640354825643807, 3.618999920488830,
    7.856013537061660, 0.9273335585580070, 2.793094514544331, 6.532912827257161,
    5.354072642139562,
  -3.273022089980290, 2.802127530707597, 5.370915950193311, 5.272385054715426,
    -1.266796131019814, 2.038632377015052, 5.865661414333271, 5.607214366019932,
    -4.745291353106295, 5.083252239126104, 5.156205293125848, 3.464494850265897,
    6.371243547375684, 3.799402329750418, 1.665328400404263, 4.076142907612085,
    2.304233683417270, -2.132692734964942, 2.185435620077936, 3.429748255092757,
    7.564117735009467, -2.458370688006768, -1.457173595520094, 1.837180516348743,
    3.386250079354908, 3.830568435474852, 6.003594742583163, -3.310648728898048,
    -0.7386163344600448, -2.223907695243580, 8.569502066062942,
    1.686286545822217, 1.315133679426281, 1.828746915630927, 3.821075853713590,
    7.704614609717948, 0.7304550847899383, 2.799569202154833, 6.457919307349694,
    5.404162713304494,
  -3.394604636474543, 2.913720635179216, 5.699800760202451, 5.000121007419672,
    -1.382372086516832, 2.001785156538162, 5.860441256288758, 5.553112253496440,
    -4.813818335023122, 5.049823398288949, 5.149415607084522, 3.227649220052215,
    6.325146767076177, 4.084391076615734, 1.263979453262441, 3.921335737365821,
    2.873637267619616, -2.089893078305054, 2.146142881369667, 3.252377555154241,
    7.854776403286749, -2.390986396958637, -1.193584883533436, 1.698774700630917,
    3.000326860187990, 3.704795878466713, 6.116441256932649, -3.275752015161472,
    -0.5261874296198512, -2.199833099780174, 8.600277436734874,
    1.741099264075640, 1.043036836764104, 1.642547982263358, 3.617899700260240,
    7.959123793839808, 1.101547397524334, 2.779066894478113, 6.547333282083667,
    4.907335002589554,
  -3.431120433367666, 2.930871339881926, 5.342557777140287, 5.591815055280846,
    -1.010139507260094, 2.117233705550506, 6.018853206373223, 5.170537020236054,
    -4.818705931442661, 5.118633922866925, 5.561068211678765, 3.266191304267365,
    6.521548195327166, 4.915115815011730, 1.450630612477745, 3.687764863340716,
    1.998095345168300, -1.905946636855265, 1.688929260134767, 2.966799053942427,
    8.517885904461403, -2.231782547879604, -0.2540578952432816, 1.405190335716778,
    2.443990213752727, 3.802640731910777, 6.102497180443599, -3.202548087906662,
    -0.3923262327741864, -1.640843278494684, 8.779797423583878,
    1.429579694786590, 1.359598030704701, 1.687564653329929, 3.343625911156366,
    8.118296761884638, 1.466688852489077, 2.467382258333610, 6.125390858438097,
    5.263008725877547,
  -3.348783268993595, 2.887160461597879, 5.564086406901208, 5.115454216832028,
    -1.319461337339617, 2.000864529986790, 5.851346004007867, 5.593461806570212,
    -4.754444800965964, 5.075374803547980, 5.234144433075847, 3.207218569249698,
    6.239160696065176, 4.025151511434869, 1.211085512461085, 3.896561557878195,
    3.041123020696415, -2.052477943050898, 2.224885088939849, 3.222005655313815,
    7.783817120634798, -2.316530131641632, -1.337176813787840, 1.793297161446530,
    3.237416178816104, 3.808643174790814, 6.010883563445160, -3.326874261022581,
    -0.5193514405936305, -2.197655376153087, 8.611995198709566, 1.727367327272447,
    1.037077928242455, 1.634513794250684, 3.629372072999514, 7.875444128734095,
    0.9739538509114180, 2.818739820243429, 6.545417859916057, 5.140073529866154,
  -3.420400029329004, 2.890461817459688, 5.590871013286024, 5.147251249987219,
    -1.264305297382275, 2.021120455622651, 6.044861131780267, 5.073527611087241,
    -4.870021722745660, 5.010092801179132, 5.526993530699301, 3.324743708391889,
    6.197456795856936, 3.846463327838476, 1.322492615386285, 3.967055946079181,
    2.928533347147842, -2.127003148667350, 2.178911411196479, 3.333811699552533,
    7.789441602179689, -2.429948889699293, -1.229535188088406, 1.661914782684412,
    2.934728403236997, 3.655027381383361, 6.160710048279458, -3.279675686304808,
    -0.5449129715885364, -2.271269846679462, 8.565515075617375,
    1.761240182445190, 1.007707396765594, 1.650377302566476, 3.664335065850231,
    7.889198659032016, 1.005162682635700, 2.773716829519737, 6.504304040102585,
    5.068924382658669,
  -3.445785492934612, 2.905440203113054, 5.864989921783404, 4.849529161542250,
    -1.625545391419790, 1.844538151765643, 5.523338742525292, 6.604553901091058,
    -3.935201609313570, 5.341714050059888, 5.188007893874851, 3.302895477257484,
    6.342287309240477, 3.980538980169040, 1.675119477810141, 4.045399723546311,
    2.245707842957132, -2.137360296552874, 2.071043228353568, 3.480732082655805,
    7.605894353769790, -2.609662109076484, -1.195829524409153, 1.685417466851320,
    3.063884474196559, 3.733776290771919, 6.060302655026113, -3.286257681154289,
    -0.5007354935386513, -2.218724672695822, 8.589027346284412,
    1.725399270880472, 0.9240552460724556, 1.589927020811672, 3.617247679547005,
    7.975988969786460, 1.203416227779998, 2.852073606649559, 6.679224830695309,
    4.586038195391292,
  -3.372090564711226, 2.899930298537690, 5.723426249820433, 4.845258835303672,
    -1.472054147970782, 1.994732335356761, 5.886734605708277, 5.606291714673612,
    -4.723929444292485, 5.097875706492229, 5.270292915983925, 3.202233557056700,
    6.246509133383948, 4.021920282555215, 1.181046784718053, 3.887550344915954,
    3.042367549776483, -2.082048932573211, 2.162538578090949, 3.100218989024276,
    7.885448801492418, -2.254207909512243, -1.269128947695177, 1.660349337350562,
    3.000643153831055, 3.745852261757425, 6.080537114779801, -3.266932766002331,
    -0.5529598013896798, -2.196293457672122, 8.672202408925040, 1.709544956389037,
    0.9777694862458538, 1.561477839597206, 3.525355565092132, 7.931793483633079,
    1.118288182789703, 2.835273142248029, 6.627958498047261, 5.020091841610141,
  -3.235050888301938, 2.919605870065626, 5.764332211767758, 4.742009974950274,
    -1.607261762530427, 2.006591715664233, 5.941311371779928, 5.699670537093112,
    -4.730810568081045, 5.145624411152399, 5.178489750423172, 3.251729796612642,
    6.404662353993142, 4.200770223180204, 1.428636849274291, 3.963431970007093,
    2.499743864483090, -2.140958738550043, 2.063623732728280, 3.444665610386801,
    7.819710779392953, -2.601913892412002, -0.9894243117926329, 1.583015374035065,
    2.787846695423809, 3.630757421991883, 6.193262537905034, -3.243703240929742,
    -0.4782879154468341, -2.187511793475486, 8.592722539150563,
    1.770338008188716, 0.9914418611478402, 1.619906891259377, 3.569460703274333,
    7.995102026798306, 1.072285012032827, 2.704770224849170, 6.500416833644841,
    5.288090769030386,
  -3.330471417610735, 2.847602002531104, 5.427890274243493, 5.276379635382032,
    -1.215063838887310, 2.009264951769839, 5.839888099947160, 5.519821666396661,
    -4.821526921635301, 5.027759570042241, 5.136473597630832, 3.427329385891058,
    6.359068008819070, 3.779580226873496, 1.506727351567556, 4.045904613366032,
    2.593113118715455, -2.131251427398329, 2.203601950769397, 3.456756564768979,
    7.611170424205192, -2.492874229680331, -1.363037377417587, 1.796239554996666,
    3.225196704449957, 3.745295073671046, 6.077657661364468, -3.297072730153301,
    -0.6582946381775842, -2.262683103232848, 8.565036163679432,
    1.735524273817418, 1.178175440859641, 1.741359163498342, 3.736780412830765,
    7.798565739490940, 0.8627850197515164, 2.787586665445509, 6.465340009952827,
    5.253878507874912,
  -3.521702132874185, 2.915659704294506, 5.564952817551420, 5.333108654879138,
    -1.114852793056512, 1.934154476696016, 5.784133047844401, 5.452210583553302,
    -4.830202471733316, 5.047299500866694, 5.125813778025766, 3.144844518593369,
    6.285735250118531, 4.100828048985007, 1.316986634066625, 3.929307845401492,
    2.895180768311507, -2.074140235822396, 2.168225765350758, 3.261778689983537,
    7.779866708726725, -2.388721539854121, -1.253431233227676, 1.736376745895531,
    3.101670981727617, 3.739440052343152, 6.071766064584750, -3.268788331437187,
    -0.6756310660814301, -2.257124966519604, 8.616193677348178, 1.689183804886514,
    1.161900262185502, 1.678479196178898, 3.618811687474263, 7.938655232403375,
    1.136886799223216, 2.760742712509855, 6.461007998679934, 4.719938334893201,
  -3.315397069861765, 2.905471420864764, 5.710962884592767, 4.897703883439262,
    -1.534354164586680, 1.970950381500565, 5.886086926207606, 5.898392529030185,
    -4.406087318108843, 5.291050248729670, 5.369205719268115, 3.012464132781460,
    6.190170933486798, 4.231531131814337, 1.172562776732665, 3.875856595205002,
    3.037710132782278, -2.055056952811164, 2.248054553939713, 3.351003889046297,
    7.699127086454472, -2.438332709951742, -1.293101047893972, 1.742524300748912,
    3.197768774287899, 3.814433894498617, 6.005159684150933, -3.300060042450249,
    -0.5347647929328023, -2.183281542773998, 8.654604970928546, 1.684901820333942,
    0.9845732445390614, 1.569523010635824, 3.530565316987004, 7.928454610344161,
    1.068703933618340, 2.803061869879579, 6.585268430982832, 5.196689243880368,
  -3.428413873133822, 2.924753496170017, 5.776463724969383, 4.945950049618581,
    -1.538639780427622, 1.837667703942709, 5.426038841826065, 6.683359251239664,
    -3.942459445042186, 5.317025039265277, 5.054172524813440, 3.129348441961623,
    6.357364767676162, 4.212968888606063, 1.366334150386159, 3.933224915612986,
    2.637516508189832, -2.067228350336679, 2.156153984096298, 3.335259522806075,
    7.661338312111529, -2.475288460467493, -1.217582343871708, 1.709481513197008,
    3.229738943189139, 3.899853719215852, 5.924751611397906, -3.297158875142622,
    -0.4343671617153445, -2.047752413622824, 8.708081211678348,
    1.721456315013860, 0.9883401097460927, 1.559193803310460, 3.519603312834311,
    7.949109100483273, 1.202905361389841, 2.931798713886974, 6.721885295365579,
    4.617589627966307,
  -3.157635423758281, 2.852289137550748, 5.591333129776991, 4.875978694336080,
    -1.462184511980174, 1.985591987350608, 6.079607275823101, 4.991080919810639,
    -5.030826370706965, 4.947505055122027, 5.185356932108296, 3.166762894120839,
    6.336136084036589, 4.309647231958904, 1.414259196121933, 3.921238591125029,
    2.587351439589217, -2.106657546399737, 2.086266195677507, 3.223253841591974,
    7.913959683747724, -2.397395879493180, -1.200479045232437, 1.709063448297853,
    2.981471467339428, 3.671880587296843, 6.141636654416368, -3.321803839361541,
    -0.3929935262345206, -2.227400397167607, 8.519914129162778,
    1.727980803063434, 0.8911189996443596, 1.612148605078618, 3.644190745107304,
    7.878255045161056, 0.8818655584442511, 2.682237718001978, 6.389706420496222,
    5.592996416700199,
  -3.394501223788650, 2.905561682912702, 5.557044894018463, 5.187466286985993,
    -1.277197998374911, 1.982019544213577, 5.729232364369778, 5.807330648139505,
    -4.694814038464802, 5.087630410534124, 5.103938245919164, 3.035115972175991,
    6.155634351695563, 4.310885695997137, 1.189054219514088, 3.816415744634340,
    3.135138171671796, -2.002991272507772, 2.185624194637047, 2.983242863319095,
    7.964120345408134, -2.154531995728944, -1.317004161314138, 1.813708561114276,
    3.243499080411703, 3.828571980411973, 6.018691369841012, -3.260363921575847,
    -0.7727097625100364, -2.168133750328080, 8.656732101208384,
    1.655021050472552, 1.365853261815563, 1.779483470173389, 3.691396814173148,
    7.848420962842905, 0.9666598436462994, 2.808800416725461, 6.527830458898676,
    4.964481577916852,
  -3.328669407784536, 2.912831215523882, 5.744323601717796, 4.822941953309043,
    -1.488923582426718, 2.012756973575722, 6.014405220646992, 5.351528808278490,
    -4.775313908149463, 5.097625913562728, 5.444946090732063, 3.294299776799704,
    6.280952088759127, 4.014027342245514, 1.324474869833967, 3.949418292607923,
    2.780528346480524, -2.109492749832754, 2.159833127171855, 3.285208719440942,
    7.814624414227109, -2.405952084363260, -1.250391551372654, 1.709052466065985,
    3.043227802186695, 3.714506838417768, 6.114942140133111, -3.264383687996252,
    -0.5222375505841508, -2.193330661915364, 8.628941966268648,
    1.759636326068829, 1.026350658773584, 1.611838591633897, 3.557559032771468,
    7.953343518954549, 1.092996441345661, 2.759778557744212, 6.548951751774713,
    5.148869456623496,
  -2.471601677080848, 2.586591829724324, 5.211026226510702, 5.056654158066756,
    -1.509273493262379, 1.893631122137543, 5.280701314498228, 6.774337589027374,
    -4.153382421437808, 5.113754823152115, 4.650175415358500, 3.073212784294582,
    6.349603279286894, 4.159632871679737, 1.197485554301292, 3.943888104832373,
    3.027236822455085, -2.051649701763472, 2.336769339275990, 3.923263252599773,
    7.239101612719496, -2.897404293434697, -1.119308590902035, 1.679981033641759,
    3.310154816018812, 4.038628253220662, 5.808867629405998, -3.407267874661099,
    -0.06325907052844223, -1.616557586381549, 8.582304039346921,
    1.355584205204751, 1.046903589122272, 1.687984505767089, 3.601137176060777,
    7.831016725038533, 0.6692157896350219, 2.452021833974662, 5.848755447357992,
    6.408077090936120,
  -3.320448388913446, 3.253709799903262, 5.172129283900001, 6.007056292392598,
    -0.2949312532926310, 1.542232758287289, 5.441676890689397, 5.730688869211345,
    -4.325302862976839, 5.373496969465860, 5.636623979811043, 3.180237678745058,
    6.160799248346132, 3.974907020735479, 1.828620235872636, 4.089226205310802,
    2.218401782898656, -2.104333113519871, 2.122740974146347, 3.431185224734256,
    7.473400102185114, -2.510877398926703, -1.318624292484754, 1.753821843381139,
    3.346402329617298, 3.914736840415729, 5.848525331839705, -3.412719583195300,
    -0.3772058474448818, -2.119513270755009, 8.504254497680746,
    1.564412201910615, 0.9205635021509984, 1.681735253783003, 3.793552750139928,
    7.733138945063793, 0.6388028769332263, 2.657692056086522, 6.133361010146085,
    5.784861638351528,
  -3.471303870804807, 2.889550773696639, 5.591758372697728, 5.187699807922024,
    -1.283263676180010, 1.975480938920721, 5.698151886733128, 5.972570081745824,
    -4.569549419266346, 5.133712040334059, 5.216426051987447, 3.265942895556164,
    6.239002103259954, 3.889461313354736, 1.196813841787918, 3.908799777380344,
    3.107729360945474, -2.060896833278658, 2.214863401113520, 3.259453214733137,
    7.766138561568332, -2.371721066685371, -1.238980292842160, 1.715059521172529,
    3.121394164562983, 3.800556446388556, 6.015835398085321, -3.304280580260342,
    -0.4877008679450449, -2.158176049414991, 8.640483950424827,
    1.711338208042477, 0.9715478659670526, 1.586366060787799, 3.587748968763533,
    7.905832167187682, 1.118948102343152, 2.889306811204311, 6.624811215325711,
    4.706152392827518,
  -3.386692958834856, 2.887901611198600, 5.495977233901991, 5.254092580031381,
    -1.202399400787882, 1.992619076557774, 5.792539195986636, 5.598641021893436,
    -4.783344424989250, 5.029693656263187, 5.204272416427583, 3.133037392542997,
    6.132656858083418, 4.057585413132411, 1.109000038319777, 3.823625804039002,
    3.319302304121747, -2.005726348169945, 2.200332541413966, 3.054576858511877,
    7.942141459791397, -2.199190008859000, -1.284202542225699, 1.791211166359566,
    3.169072642920213, 3.792392662590062, 6.036041633770368, -3.328394251003055,
    -0.5415256528478126, -2.189783019703794, 8.605194447746470,
    1.718124418154977, 1.110139045222000, 1.681600256712513, 3.663549782872161,
    7.874047671158085, 0.9838146905142050, 2.798314767207644, 6.499834182655383,
    5.057281871916913,
  -3.268373847640958, 2.775665019996381, 4.930030065862932, 5.786709482990446,
    -0.8207035001165758, 1.883672790713845, 5.554579365520583, 5.995034224927066,
    -4.593474600804331, 5.086092216404198, 5.129371789409306, 3.280609705564465,
    6.121050718296882, 3.687346678404643, 1.325873360326498, 3.937138061408690,
    3.220689358989527, -2.087798057827904, 2.224991846233522, 3.064792526893013,
    7.845760743129590, -2.265032153005679, -1.496551195993952, 1.740538203128099,
    3.253194827490010, 3.894684805550730, 6.313363849150164, -2.741931395532526,
    -1.353485359836765, -1.214764098872883, 8.785354681167092,
    0.9343015266555156, 2.370075867832242, 2.249739622028697, 3.616824141944588,
    7.679493200758508, 0.9180439110761311, 2.663051253954738, 6.132015303507264,
    5.694853961279568,
  -3.427453923566583, 2.908947284265641, 5.350641787095170, 5.662067627303108,
    -0.9135710838296526, 1.332020956938583, 4.957064323246763, 7.023918527785743,
    -3.293829971332641, 5.630657111771455, 4.757001646571512, 2.130909052522952,
    5.937913928690900, 5.423821610832465, 1.037153476408099, 3.637554191892938,
    3.159914944711927, -2.001842484044265, 2.008164111304514, 2.631468537999505,
    8.411002238883718, -1.878545102468967, -1.119528714480424, 1.702594209173103,
    2.822825654818391, 3.634855728282775, 6.211456475971474, -3.212801843122296,
    -0.4383162911139465, -2.013367235228874, 8.601200302343873,
    1.794009517475585, 1.176871560655322, 1.748671540928034, 3.662871340349837,
    8.016002936377147, 1.318301229335681, 2.761479569984862, 6.362226482512108,
    4.336651911304727,
  -3.337659364690654, 2.906068788333424, 5.711958822882010, 4.913808454681599,
    -1.527508581384799, 2.005462184802248, 5.957393624762719, 5.765679304425273,
    -4.448627487222191, 5.279532052652636, 5.454819459284606, 3.118216865308221,
    6.244999554203296, 4.225043947186795, 1.300352256337293, 3.912572347555255,
    2.769024766330525, -2.090142707786063, 2.176781933559891, 3.317317181564400,
    7.783532295745991, -2.436590761971768, -1.266410329678103, 1.733970556597950,
    3.108690522377325, 3.741075927973236, 6.085324724761713, -3.273367154807858,
    -0.5720564167485384, -2.222152863102654, 8.631456695838711,
    1.751618340056111, 1.050448896549998, 1.621179941150318, 3.576462083793211,
    7.917511398970261, 1.044181453699214, 2.785872998898336, 6.567700714016457,
    5.180606587536719,
  -3.425746942037036, 2.903836673930281, 5.606822394848761, 5.156752289639901,
    -1.349272354320984, 1.987438289228610, 5.763534954508409, 5.999464017803310,
    -4.494328645991121, 5.202557005423987, 5.255157301030768, 3.201186957332256,
    6.259278537320033, 4.010418404764817, 1.231022896620221, 3.923942438794893,
    2.984781207639722, -2.077533913554619, 2.216441632859703, 3.363672600998814,
    7.738057583430301, -2.454835959762918, -1.230841880735396, 1.736446786765073,
    3.114561465251882, 3.758241800667542, 6.059998925673073, -3.305529872041065,
    -0.5140708386343065, -2.199668875853536, 8.593107522823797, 1.747651631009713,
    1.025952612693553, 1.648386018405113, 3.665566558348176, 7.886105831370116,
    1.021824365923348, 2.846287501051537, 6.591243383317622, 4.873250075985949,
  -3.405748942545659, 2.899080093369625, 5.604815394657217, 5.118936340650281,
    -1.350575637996021, 2.006254117956864, 5.831181363982013, 5.776464815821471,
    -4.628022999034804, 5.153476708599365, 5.250552146120503, 3.180222159062879,
    6.262810504949683, 4.096681539634633, 1.231423636522762, 3.899878094336479,
    2.945862274609507, -2.072258271774877, 2.180349367468104, 3.162920614396740,
    7.865834026112676, -2.295050973965115, -1.297299288061857, 1.757755565258625,
    3.130513537945166, 3.753328660822357, 6.068900028317518, -3.292438956985383,
    -0.5898544698166650, -2.235117797902388, 8.611754517283716,
    1.761067422211268, 1.086188620766420, 1.663506805310983, 3.662872895594738,
    7.859045160216522, 0.9801085115007692, 2.850929031481167, 6.595529852186818,
    4.968249404432111,
  -3.363608943894988, 2.910344299240985, 5.737616367916913, 4.868343022285480,
    -1.475160511034364, 2.021120142049722, 6.026408116995113, 5.398582021992010,
    -4.698192583333918, 5.136641599429608, 5.532981951509903, 3.297813504206496,
    6.237994811452290, 3.946287453912805, 1.317828952022751, 3.952375407117378,
    2.839275522666712, -2.114854852124630, 2.147124242531510, 3.215398685076403,
    7.863358472990040, -2.353897337891592, -1.237415013517166, 1.673121738642469,
    2.980470256956500, 3.700519180162073, 6.127644031356901, -3.255550523508806,
    -0.5592053948971011, -2.215489662057907, 8.634129777107983,
    1.771058902452621, 1.055904898325135, 1.626068266804784, 3.569520736885068,
    7.948517073081726, 1.099690555043747, 2.769105112056785, 6.558838707013090,
    5.095883458060640,
  -3.357024545322157, 2.901476775677018, 5.717305861293503, 4.844694895842595,
    -1.466954735179449, 1.981495256819056, 5.864150397084424, 5.628867940001839,
    -4.712018228431264, 5.086040574173441, 5.253044853294588, 3.089038510424260,
    6.131099119853067, 4.083641646154525, 1.090496420572943, 3.810250476367249,
    3.274272370107838, -2.021334974919331, 2.177598212595992, 2.915535298872271,
    7.916293513003835, -2.094390865739962, -1.358789760633664, 1.713377971311943,
    3.140149671063969, 3.835844665052925, 5.982588570153232, -3.308558659385000,
    -0.5408395817384749, -2.158374805403302, 8.683736934674995, 1.597254629132851,
    0.9377041848611967, 1.529063138536486, 3.519632288619035, 7.918036086489477,
    1.092642313003589, 2.851912793871833, 6.644005546806174, 5.053840881453556,
  -3.305146837250507, 2.905588573921460, 5.690081914003835, 4.677994127551513,
    -1.464906929401315, 1.933943187733909, 5.328215181406086, 5.728781373572872,
    -4.646215809424976, 4.671721532290633, 3.964216141468054, 2.168071589404197,
    5.665512640659586, 5.083909353140508, 1.078040717935343, 3.653058705416274,
    3.744278559634156, -1.921835588174674, 2.061409370287823, 2.937974628727935,
    8.633367006940194, -2.035590137787896, -0.5140189958008424, 1.782618352884436,
    2.746385321008853, 3.728847884016869, 6.139737035499891, -3.327073457533950,
    -0.1775671277938340, -1.839942229463185, 8.639000632458652,
    1.516646782438226, 0.8388426033087849, 1.532813480763665, 3.549920840171020,
    7.931704128165860, 1.034438393776729, 2.802768054558205, 6.598563769186975,
    5.149388431465654,
  -3.293725500947992, 2.915034094311107, 5.760611705628740, 4.743450919993967,
    -1.484044623732061, 1.962341708995493, 6.047937533895770, 4.987532115466962,
    -5.001257064867529, 4.946754712649999, 5.243982454971094, 3.263327808530487,
    6.389745214735895, 4.153957212142957, 1.380911554633392, 3.971078104924023,
    2.594203650770002, -2.120441633012763, 2.184080475410834, 3.612357554081627,
    7.553725614455385, -2.661830204959291, -1.206210919428108, 1.705507418659535,
    3.122587521112008, 3.786438189536002, 6.060114107816350, -3.304733443959680,
    -0.2870614866796306, -2.010748120703881, 8.616176767880397, 1.668736388161801,
    0.8760924172323655, 1.558880493899100, 3.530174772229578, 7.973324749497666,
    1.104525212051058, 2.720591294513231, 6.509368711648039, 5.266871132631616,
  -3.449121860251388, 2.937771192052196, 5.690121415899738, 5.059167753516063,
    -1.313919430499290, 1.956109065168067, 5.952142322563967, 5.186165709167890,
    -4.912254447596425, 5.032073090628405, 5.127940920584551, 3.120651162057083,
    6.389552725065709, 4.296140567255315, 1.404812643555836, 3.939761575805407,
    2.557063031190931, -2.106612068025762, 2.093471631325056, 3.294416237130213,
    7.810313239410458, -2.442618417657999, -1.206930486942763, 1.692944258400511,
    2.987498261941801, 3.670872323991860, 6.142468938784408, -3.266450668813913,
    -0.5904761453258918, -2.280666565360709, 8.582516952338962,
    1.784928943171605, 1.061450685424879, 1.659218188246554, 3.646825179222699,
    7.903250090409985, 1.015024271843123, 2.773828390651305, 6.525810663791452,
    4.991474666396181,
  -2.549913271865330, 2.514755203794770, 5.225908284766071, 5.165718851589875,
    -1.563491217121799, 1.955099476034174, 5.810630810784284, 6.124720897052144,
    -4.144922300887528, 5.426376575349559, 5.320315908518755, 3.115097822368061,
    6.373886658164905, 4.587892706101954, 1.743642974253766, 3.859446737014274,
    1.931157580691571, -2.086473550505592, 1.815584672103406, 2.514746964129301,
    8.357491237116768, -1.906467675238027, -1.279383731287879, 1.610708024523446,
    2.734973124445293, 3.523516868756284, 6.237880557543416, -3.212456473708384,
    -0.6859173593570688, -2.438843361719182, 8.525074225084783,
    1.797457836652606, 1.094064822257917, 1.667126502660429, 3.579560166904993,
    7.652515635425569, 0.5903467576234770, 2.519876879114698, 5.883523457705547,
    6.496796939127987,
  -3.443067406569380, 2.902015911547958, 5.656828810579785, 5.073384994739182,
    -1.472724151380105, 1.960598982283709, 5.557950547795338, 6.507127957861583,
    -4.043516470270123, 5.266541149949219, 5.143727510831664, 3.478859446598432,
    6.382770560488697, 3.868163985388686, 1.829374562045658, 4.052186664413834,
    1.920028389911435, -2.117005185474952, 2.101858230934544, 3.113489645573649,
    7.617568904484258, -2.192580048708455, -1.625247969748007, 1.834809911775006,
    3.537184388521252, 3.955374386866523, 5.828771682496189, -3.370935680781906,
    -0.6104997263775506, -2.141401185731672, 8.550094919514862,
    1.628815170637263, 1.236632167027665, 1.827834989531207, 3.925557897801477,
    7.753098117659183, 0.8058700854860640, 2.858089905921330, 6.639511875236638,
    4.778236932843739,
  -3.324429177553240, 2.887228740854793, 5.625386268578846, 5.024343298961830,
    -1.443004462162716, 2.021329127221937, 6.009737603290358, 5.552508091291465,
    -4.569191864866432, 5.221653218308813, 5.506755617522427, 3.123657777951617,
    6.193210150162151, 4.150201529772919, 1.266871340772016, 3.910241688685238,
    2.908565451505243, -2.065182273085838, 2.224704033530087, 3.361697884591383,
    7.713708589164450, -2.452787993951433, -1.292476789442493, 1.764348188374530,
    3.212283112201432, 3.807057803624193, 6.016654307411276, -3.310037890216374,
    -0.5647679819557445, -2.208101003162488, 8.638493618565581,
    1.661754567634145, 1.030054580543682, 1.595759126540324, 3.548219187896686,
    7.919158518370292, 1.052205016882470, 2.760772625537300, 6.507646863861964,
    5.274042426481499,
  -2.658711662783392, 2.660494456563432, 5.281491052227752, 5.129334459316290,
    -1.442731054188984, 1.902483679046335, 5.676713220074196, 6.260676576628184,
    -4.291349182164173, 5.283219181520884, 5.261416262706033, 3.297218773057658,
    6.235591056186263, 3.664680740411380, 1.369776722275500, 3.950955042061028,
    3.150660418030319, -2.095155870624376, 1.669036459983971, 1.829365187534377,
    8.904324196756567, -1.197013544213871, -0.9452909912446797, 1.509915988614309,
    2.394202249185998, 3.461233299594346, 6.293667786440843, -3.172026339014605,
    -0.8086303293789120, -2.450392930187117, 8.608192963298263,
    1.746883158554747, 1.144858305918080, 1.628621299913623, 3.485899166616746,
    7.792352862316020, 0.7628665981390786, 2.564693464954871, 6.014866086452314,
    6.315336900626368,
  -3.432302287910984, 2.462530832947668, 2.842651588594430, 7.123080063665865,
    1.198914235051517, 1.425394525483508, 5.116925386834650, 6.116824244811786,
    -4.258230977081794, 5.309063034589635, 5.474272489481283, 3.183482862339595,
    6.330024289236543, 4.266070613908673, 1.244439108546594, 3.889254459492454,
    2.795665432386329, -2.122252376594676, 1.916093374363329, 2.442246336213360,
    8.538307417025113, -1.683188078236379, -1.188477084885517, 1.681496626736752,
    2.685835627593216, 3.525549829836285, 6.306330284328022, -3.236232369153042,
    -0.4148706920212273, -2.007715289651423, 8.455492391172813,
    1.710819972989910, 1.090048798383633, 1.843764587737005, 3.830194444549447,
    7.484488961479705, 0.3491353382948571, 2.730616734617477, 5.453435200830894,
    6.122790904772224,
  -3.264718738331240, 2.883462726762825, 5.562505693328351, 5.031107504662857,
    -1.412718046723834, 1.972245782170611, 5.740226797371873, 6.013609364473039,
    -4.521669624043227, 5.169054264131120, 5.197021576868674, 3.208574026196576,
    6.233411301687005, 3.946804823870812, 1.217436356001639, 3.913442741157764,
    3.077065302016561, -2.064410487341748, 2.224751814096526, 3.281157619915090,
    7.748309482880063, -2.391477801462460, -1.258711521683575, 1.718817914014771,
    3.131928942732649, 3.790098510857280, 6.032647572250688, -3.283027965872654,
    -0.6091597764905030, -2.233510169940871, 8.668659403151523,
    1.715711675343316, 1.052892526982732, 1.587783201818966, 3.508294751727603,
    7.919532299589827, 1.065781064720133, 2.784616747501604, 6.510786475773704,
    5.304674408797013,
  -3.370965190402948, 2.912279435913534, 5.751453314407105, 4.848753064391234,
    -1.453133856559407, 2.024346146440195, 5.903646797139997, 5.598280780970712,
    -4.607084619334601, 5.126135910969054, 5.490304266058684, 3.380711318654416,
    6.261339142598513, 3.787836303769289, 1.167168050008368, 3.924487030051759,
    3.024898209110869, -2.082807048429946, 2.197390519849958, 3.038086533255339,
    7.938023268630898, -2.137822706277794, -1.424532418376803, 1.838310909523321,
    3.248655665131979, 3.795511207623942, 6.051627584755590, -3.338374613928026,
    -0.5095517976194993, -2.169571564877860, 8.603087733811495, 1.781531423613349,
    1.139093994144990, 1.715896179454820, 3.735684973370296, 7.831775473919124,
    0.9252626848308531, 2.855859119717532, 6.658117306977354, 4.957641897069865,
  -3.200903882888889, 2.987780965951991, 5.135794017848763, 5.736082309174707,
    -0.7572896421538601, 1.836612859596803, 5.557066471388161, 5.568232559656954,
    -4.469240183851293, 5.304614757790993, 5.155219298431018, 2.393541920821365,
    5.922405235187125, 5.376653195987819, 1.461540308838479, 3.761840738699401,
    2.311687518911588, -2.044275869309235, 1.914467230950390, 5.412597387658604,
    6.032104279804201, -4.142963750333727, 1.125802879294512, 1.788112647571359,
    2.202418449596630, 3.385519393522211, 6.394382544899226, -3.032138615661640,
    -0.9863651672963929, -2.269877883671586, 8.636751142766595, 1.656851217035626,
    1.409286312874167, 1.786470019046106, 3.631840862372308, 7.750516445087994,
    0.8209242386466892, 2.683631615574532, 6.189346457037072, 5.863493567553899,
  -3.581429275947816, 2.773768591976700, 5.734748585331443, 5.024794135055004,
    -1.428342645295168, 1.972531490680920, 5.640934023960982, 5.959930765212632,
    -4.721131484013242, 5.014462222303200, 4.717821446031008, 3.110535234396780,
    6.458171413120515, 4.253365020080210, 1.223851647546461, 3.913040997163225,
    2.775690476052143, -2.056933727439459, 2.168897174333782, 3.456279262157354,
    7.633284793610271, -2.559167735317606, -1.149043483239895, 1.713318354032242,
    3.120788776440494, 3.799155427495698, 6.003222307460261, -3.309391882425369,
    -0.5372118829465845, -2.192229193890447, 8.627685758735574,
    1.616921079588120, 0.8988210783150912, 1.547818678718627, 3.654405781320442,
    7.843184605008823, 1.117555273640021, 3.011910867554639, 6.766605096857737,
    4.026185802363495,
  -3.414779152833816, 2.894976187936974, 5.570528521637665, 5.166677016683772,
    -1.307480479241294, 1.983855865183004, 5.749467834888443, 5.949623002765844,
    -4.546191630493256, 5.159008716026290, 5.287248116524057, 3.236150681284015,
    6.191905638053123, 3.862434804195031, 1.159236165085454, 3.899711238097753,
    3.211159194872835, -2.066789208050971, 2.233298680451051, 3.302959233550744,
    7.782601547184100, -2.401786767358654, -1.227263452276563, 1.711559099818225,
    3.056043560527967, 3.736118988647527, 6.079193701679979, -3.297172182609692,
    -0.5234728510578213, -2.218326506017778, 8.600658325731477,
    1.740269984465318, 1.000910849564383, 1.624827751424342, 3.630096649433058,
    7.891047491720245, 1.050103845273300, 2.837077063426512, 6.572929745261549,
    4.926872685332206,
  -3.406481680405466, 2.960285657240808, 5.762311295377669, 4.997775636920243,
    -1.260441623990817, 1.904672182938085, 5.725335544366203, 5.393934261215182,
    -4.883076392653244, 4.954374144622914, 5.027118593100822, 3.134984847804098,
    6.240620050104908, 4.114762019139237, 1.279380153582595, 3.887719205175713,
    3.016323372186049, -2.090057422401703, 2.116862090362106, 3.052505917678878,
    7.928537974430488, -2.242843602509938, -1.259225137987848, 1.628391320478083,
    2.882836514902573, 3.640093270125301, 6.175331878176736, -3.124636552725752,
    -0.9181960630724371, -2.251675061918829, 8.694273935264681,
    1.588959656790218, 1.359659236581529, 1.696009661025925, 3.497661798683489,
    8.035765137313497, 1.326465130690597, 2.659345903114542, 6.418776459411405,
    4.816881864344467,
  -3.321050155728335, 2.896764031481006, 5.672013259800779, 4.905218069631987,
    -1.414957541901651, 1.992387173206247, 5.916163181669424, 5.415213050278277,
    -4.827749337836677, 5.036166758443389, 5.281928851742634, 3.271268631962319,
    6.257729644925832, 3.948466922295166, 1.246196809428332, 3.921892396168029,
    2.982563398469452, -2.079723341763897, 2.201142098078815, 3.243951024684932,
    7.772445229582035, -2.347199115746123, -1.295775609053235, 1.718701640841596,
    3.122501218268225, 3.783912345702086, 6.041923455068835, -3.303324445550015,
    -0.4713546338358643, -2.165368908339254, 8.636722535489509,
    1.741130778414773, 0.9833815763731590, 1.593283362971014, 3.562287168076317,
    7.930803814945777, 1.057224276447692, 2.794396636355693, 6.560689516541077,
    5.168756690698754,
  -3.242398158303248, 2.736598264932288, 4.984724054733660, 5.652873005323381,
    -0.9886845973622606, 1.984079994438830, 5.476103657412497, 6.264963728331271,
    -4.499940005389100, 5.060097614465364, 4.960746619818026, 3.422410380318288,
    6.365220909569279, 3.755119974794733, 1.275514680970905, 3.944857235701849,
    2.949716376281021, -2.152759225352142, 1.990009502482414, 2.644273005516026,
    8.304445939974450, -1.898632132785871, -1.194070950876942, 1.576745763159509,
    2.669564373445614, 3.545924511326492, 6.260393304065349, -3.220019815072662,
    -0.7361577079299252, -2.374413021435079, 8.582155811265277,
    1.880904895812741, 1.197536517107079, 1.745676275914032, 3.668645794043057,
    7.732745296654251, 0.8294029966922745, 2.764181761153112, 6.282821065971136,
    5.597888588776123,
  -3.026058910231666, 2.802928172681041, 5.475986352761138, 4.958367683930407,
    -1.517502428781647, 2.043827693585257, 5.912265861772640, 5.850331515292291,
    -4.476640404926647, 5.233113040573458, 5.319581798026584, 3.370340695032631,
    6.437662592903542, 4.151433774516979, 1.574575726361586, 3.958953495513603,
    2.099495542071660, -2.086234633070729, 2.036149960555474, 3.384796601789165,
    7.619118490062815, -2.524907082360459, -1.271165337290372, 1.642688029761530,
    3.060970169181491, 3.782265871672374, 6.068301437416236, -3.235215376169688,
    -0.5983886589791920, -2.061732198250625, 8.679859658533806,
    1.667553457739788, 1.189118456341022, 1.671915849108118, 3.509202264918365,
    7.937946425618102, 0.9374078732048399, 2.621302808708636, 6.262379720215534,
    5.872915022563245,
  -3.293013214937258, 2.879109224557403, 5.592120786454227, 5.011320798630336,
    -1.419322907602842, 2.009837067009022, 5.906895971231273, 5.641424609673419,
    -4.674514941808165, 5.141688269859428, 5.293277921914300, 3.145247277233123,
    6.231228890640176, 4.119138594203133, 1.203070922206507, 3.889908750750004,
    3.002165544032870, -2.058068506357383, 2.230767577518008, 3.247085834226788,
    7.778648988641862, -2.337159999883539, -1.349737497343387, 1.796164011272839,
    3.238903748324147, 3.798073943074106, 6.024556009765784, -3.321328524901217,
    -0.5535065689980915, -2.223873305248336, 8.611899374389047,
    1.739616498741634, 1.060585177247194, 1.644854328447405, 3.633857610833523,
    7.856764608944039, 0.9341261950728575, 2.803223397159302, 6.539573495923611,
    5.276171246585322,
  -3.264389309715101, 2.882055320653205, 5.534853865739928, 5.089051276266695,
    -1.302745772094184, 2.011206802751391, 6.154430441769760, 4.724796101227150,
    -4.953327593328450, 4.919526940854207, 5.538600248372747, 3.054498264673003,
    6.102775390382526, 4.287990372657619, 1.169896387254792, 3.826033734669632,
    3.119276084091556, -2.063371462818486, 2.096283152558794, 2.817288624458239,
    8.179025327579801, -2.024760121329259, -1.306564289983531, 1.748990733294288,
    2.977174238247198, 3.666923136888356, 6.158590671175729, -3.314974861944366,
    -0.4694133975880816, -2.251487311106676, 8.558710337493567,
    1.736561536975790, 0.9959221905898670, 1.637168133479224, 3.614687043026963,
    7.879981077593249, 0.9501205934527928, 2.659830856757192, 6.343371674098806,
    5.506208758763153,
  -3.228261960662735, 2.764842750252672, 5.134983351996978, 5.477678653679686,
    -1.232699695880306, 1.869802096089344, 5.146349539743797, 6.940273797677880,
    -4.068417256128802, 5.061063126700802, 4.628345855843320, 3.381705443714196,
    6.463633136419769, 3.742142775692220, 1.450986434333837, 4.084081058900532,
    2.662335550146666, -2.152847883163085, 2.233678693095687, 3.927705986000320,
    7.338696574849235, -2.859430229715167, -1.129751849148931, 1.729902255390108,
    3.047018203248871, 3.677657449978038, 6.149988183280148, -3.360927619141928,
    -0.4045441290719534, -2.247901700124441, 8.450347484484579,
    1.799347291689892, 0.9547843105229517, 1.719875239533666, 3.869860913499232,
    7.643158794689069, 0.6453959864506149, 2.890369721436359, 6.483428602742773,
    5.331397973331074,
  -3.363076212158083, 2.913720156318670, 5.763301087930388, 4.820560478758499,
    -1.570475435293337, 1.987996157454945, 5.767771380094472, 6.075415968162017,
    -4.423517359307290, 5.225512806476289, 5.185720976220729, 3.329897460098053,
    6.377971051559831, 4.034954681366425, 1.546047825314482, 3.982667154620784,
    2.386719387260968, -2.105611609048517, 2.048434188099017, 3.049075867935365,
    7.881094441729576, -2.255424245107746, -1.299242698588774, 1.692604534020476,
    3.069165986963963, 3.750575496422604, 6.071449521369344, -3.248485359573096,
    -0.6939976773734314, -2.286177283366889, 8.674258113752398, 1.785866988881071,
    1.104517433008094, 1.625043855511619, 3.602472549665574, 7.861584581339306,
    1.004975483832427, 2.903500654818452, 6.711228951707869, 4.966895241756079,
  -3.113111561940883, 2.809075271520434, 4.110757284081719, 6.633796128038629,
    0.1859638829994180, 1.601681493988317, 5.335912610991926, 5.853531367815411,
    -4.576411900619280, 5.215109348099213, 5.093182994260590, 3.095543019562578,
    6.436721806523678, 4.225931741374541, 1.335591224030240, 3.907343254257545,
    2.555522244377916, -2.130279235780038, 2.180642703057718, 3.031324359870756,
    7.700449053392723, -1.875735965769526, -1.961681936770394, 2.025570208225074,
    3.669693068424065, 3.963770863291045, 5.843956822218393, -3.461203348732120,
    0.1346065351995216, -1.425535468911914, 8.386105262535455,
    0.6525874462993522, 0.5558752132505641, 1.537472382952536, 3.702469099093484,
    7.702191919228118, 0.5551723220240345, 2.289638908898449, 5.335544729096878,
    6.370529606222863,
  -3.316114769393852, 2.896126316649937, 5.658410860137630, 4.926579667344995,
    -1.394129559902938, 1.986163054077597, 5.911635215934660, 5.358834501058314,
    -4.866175521062097, 5.009500028477854, 5.242242813346691, 3.262313981796221,
    6.272528794755742, 3.992114591660396, 1.260711862577519, 3.920187352067376,
    2.945441120239813, -2.074636684255432, 2.210241639912497, 3.241507455768695,
    7.759547985830864, -2.330338950983295, -1.345784200505737, 1.769479486925524,
    3.207269311444137, 3.799612019103763, 6.021649778567217, -3.321043032496127,
    -0.4444770583939017, -2.161852372758918, 8.619411791308410, 1.732762856553396,
    0.9599430056153473, 1.591677849105432, 3.581124886410500, 7.912930897425618,
    1.020886463002318, 2.798736358323636, 6.557302971891874, 5.190332586511742,
  -3.638743046190718, 3.107163237638625, 5.114297016491928, 6.018619749427218,
    -0.3202829750647330, 1.664433205182572, 5.312605492799582, 6.029489454347466,
    -4.232024844016427, 5.262401797713435, 5.614171430044214, 3.672115941515768,
    6.335493977821586, 3.858879378217768, 2.009647633956387, 4.049219554263036,
    1.627149049653046, -2.088144771137335, 1.920614228566192, 3.424321826535911,
    7.570333045452858, -2.558983896024754, -1.293101774718884, 1.716257334472009,
    3.127215700457105, 3.764570117574435, 6.075352305375522, -3.284855174208899,
    -0.4574363827529273, -2.039465351247935, 8.580777077685612,
    1.579622032257248, 1.118113177407744, 1.683982426157812, 3.586265683160537,
    8.067275773881404, 1.214442058674500, 2.585470300767918, 6.115632733291362,
    4.611750625405286,
  -3.485822282493056, 2.913619896205773, 5.508631150738180, 5.274946845879010,
    -1.187551786808023, 1.921717817926579, 5.795675158360917, 5.531432851032640,
    -4.752237904597625, 5.110467302820383, 5.031319598546387, 3.013250852868895,
    6.316684683790960, 4.271491945679428, 1.361892847679273, 3.933679215494996,
    2.737308483669708, -2.108054246670452, 2.195795861936423, 3.160925541204464,
    7.744546690611385, -2.312870203380773, -1.476825853103754, 1.718093360104207,
    3.278409772568316, 3.926070389226055, 6.186113967352139, -2.941431222447731,
    -1.203803452939931, -1.478077381850888, 8.728948860296798, 1.201183328696766,
    2.145072702055167, 2.275262341201222, 3.910025800863109, 7.579372350414928,
    0.7460248080314190, 2.844187096086888, 6.544065701309528, 5.014748434347437,
  -3.368313326434238, 2.845156520634931, 4.857170594529003, 5.967390624427335,
    -0.5634732658251178, 1.787250983276444, 5.527136714678247, 5.548157453523477,
    -4.782625720315012, 5.014639317600846, 4.898829854435608, 2.608592974095908,
    5.910721875270249, 4.624146069125264, 1.080929835892675, 3.675965259388661,
    3.530672847203021, -1.893502978166775, 2.281343174685643, 2.892743207256720,
    7.813641689068037, -1.934640270181616, -1.645602751259581, 2.018692179040874,
    3.756440329095617, 4.036572219225983, 5.712436316601795, -3.538823928093004,
    -0.2889138273335403, -2.082336415605049, 8.497322637082730, 1.446109975731103,
    0.9121285400629042, 1.656000093913541, 3.798930271912849, 7.639786347132148,
    0.5825465573902906, 2.711644701651310, 6.134586903453359, 5.728612966117026,
  -3.016108021108444, 2.812229217599487, 5.656930723222164, 5.069791868766849,
    -1.548666137236980, 1.745630353644367, 5.851607134676438, 6.015838304740440,
    -4.122040057103064, 5.583821425568477, 5.179390264931776, 2.083221122536114,
    5.734263616173410, 5.039045037608337, 0.9611143734093692, 3.680006405289621,
    3.755272961765608, -1.841067916501273, 2.423197606040130, 3.742525829950980,
    7.421568082626582, -2.780680283706324, -1.076569184724758, 1.779746134628765,
    3.410194197640239, 4.028224299386473, 5.777948982763793, -3.417094241036715,
    -0.3341424688295063, -1.972632607543752, 8.635959538120888,
    1.471837979145412, 1.001357637099292, 1.590745035298455, 3.483712612086884,
    8.004965249260701, 1.053397443185166, 2.551532971189555, 6.269191523654727,
    5.782918610086351,
  -3.318687538286622, 2.867242874619827, 5.592068019063230, 4.972193739807536,
    -1.414242983959388, 1.976869358965733, 5.834478879404456, 5.661722704277806,
    -4.763798534028982, 5.068783351298523, 5.116278288159546, 3.231212875194961,
    6.282002198848144, 3.984885728470362, 1.329198910834968, 3.931743946246190,
    2.861206107418157, -2.089141682926380, 2.105703839873350, 3.061373002339759,
    7.877372758479500, -2.281400287444341, -1.196812859483524, 1.599974357632034,
    2.937658060818896, 3.756470205660108, 6.058267538383094, -3.242168093359533,
    -0.7250990187836471, -2.260020283151451, 8.717590036738020,
    1.511125591115082, 0.9440066536470221, 1.479705078444835, 3.423995620141369,
    7.925194295880727, 1.150688481652044, 2.816104791534927, 6.561885211883504,
    5.226213024880483,
  -2.844195814022281, 2.724854943686345, 5.312147870023384, 5.129142066746695,
    -1.425861202493095, 1.924090603998389, 5.639986932097639, 6.335466983565859,
    -4.321810808738713, 5.206437089675574, 5.171050733252839, 3.423578086579143,
    6.237696400147652, 3.576187172759250, 1.560137225656136, 4.106395270371758,
    2.732590881358027, -2.134155954452070, 2.198484534508437, 3.705504400990680,
    7.437921143570546, -2.788538099853214, -0.9894913673343747,
    1.552377025222869, 2.944314115991364, 3.813474778461121, 6.029389304187044,
    -3.279688648170207, -0.6071965317850296, -2.185279664819796, 8.713638983488492,
    1.594647599094584, 1.076782061989235, 1.536905653484679, 3.296680769541968,
    7.971432166306588, 1.085493473628899, 2.521438108024108, 6.067705202926910,
    6.115026312258587,
  -3.555575456596137, 2.911771698283906, 5.476713065546729, 5.533129723070452,
    -1.000805394726952, 2.016094874090165, 5.927336541915432, 5.409005701411594,
    -4.621274387100028, 5.092688821174356, 5.974388957208063, 3.980044718201203,
    5.492351798358076, 2.947658578490461, 2.635730115788707, 4.556935280474185,
    1.764023843652530, -2.169828384687185, 2.050216600983398, 3.609743898481475,
    7.563329122984608, -2.821078748718519, -0.6617085170995222, 1.720192389210196,
    3.403683861975818, 4.257679225831572, 5.524553666603604, -3.483097917274551,
    -0.3333177570710101, -1.758455740119371, 8.690907080437761, 1.147687693442956,
    0.9444978273715007, 1.524108943570588, 3.532816002825106, 7.984444049785986,
    1.162582431779388, 2.797248407660281, 6.475370770990306, 4.825759190619126,
  -3.474025894467327, 2.905251941495852, 5.732205250477114, 5.038578459129075,
    -1.458622650762214, 1.873618359372932, 5.458371913174728, 6.607397438909969,
    -4.072750161810965, 5.260592861867153, 5.078670345271678, 3.250897175666135,
    6.331276950208288, 3.946624454702818, 1.384539802729958, 3.978094760808075,
    2.742287485268349, -2.094575516032767, 2.152036736413356, 3.285635498907125,
    7.736092818081080, -2.422945382253198, -1.233797438108224, 1.722892193483020,
    3.138439007518078, 3.791614731806978, 6.010494349518707, -3.295023008316451,
    -0.5270676662891950, -2.195407817455224, 8.627336892450561,
    1.741447953149164, 1.013779292317025, 1.614016768298302, 3.614724477306910,
    7.939351617744874, 1.202305059884511, 2.890518466722777, 6.655928475786270,
    4.450629353006457,
  -3.161390482688333, 2.820218753835406, 5.503957117406767, 4.959470759473421,
    -1.479851381216351, 2.014781023888230, 5.812340895048719, 5.818777727839945,
    -4.780063937522649, 5.050855699939918, 4.987295921792956, 2.693538805322783,
    5.898337267636027, 4.987126463807943, 1.299871922227103, 3.678406301302007,
    3.169861192787534, -1.968025814199265, 2.097192973835061, 2.855217597241803,
    8.338682844185799, -2.080487275368633, -1.000656705948591, 1.769986691202491,
    2.958776248768593, 3.715100038847866, 6.076562353422747, -3.345145135833799,
    -0.4070570654973968, -2.183799732916381, 8.495375776437994,
    1.749621641188894, 0.9971181437325054, 1.727384309665400, 3.848502934147322,
    7.712057301322033, 0.6412077718997249, 2.781759515914713, 6.480356593258489,
    5.493502373870428,
  -3.412184591787371, 2.899312801682036, 5.675887807788005, 5.031951001056434,
    -1.425301948972345, 2.018714890761380, 5.847233233780504, 5.774242995906579,
    -4.650823779018927, 5.151820214860072, 5.189863084983265, 3.239722400711210,
    6.347975165427963, 4.095021545950703, 1.346326093813074, 3.945734182705085,
    2.691215897183965, -2.082646650409560, 2.175726366512087, 3.355582001538086,
    7.703548589081097, -2.455696760028744, -1.282605528743817, 1.767539174470240,
    3.209641771036738, 3.799818918596694, 6.008988616239658, -3.332613118792104,
    -0.4537366768871722, -2.178467255052017, 8.583684126782483,
    1.717012199453442, 0.9587179301513954, 1.618870777966252, 3.659585887545667,
    7.897820819259708, 1.022666460637550, 2.840459883200239, 6.611535720933438,
    4.898503355142389,
  -3.619799089872022, 3.085797033948352, 5.961796693836493, 4.907543410604538,
    -1.446129641183646, 1.694237527445268, 5.562234588865881, 6.012887071706987,
    -4.593234029007585, 5.229237535139065, 4.333570288480406, 2.357052443090456,
    6.382298758587130, 5.461390449397793, 1.385641087831014, 3.715526138721827,
    2.214502669081452, -2.036925589535504, 2.007106606340005, 3.635984078153039,
    7.507623062314882, -2.843856536086367, -0.7602820712174366,
    1.450029720455133, 2.814033460393405, 3.860884032784920, 5.993705038942163,
    -3.234575987815894, -0.4980338273778442, -1.947205035461523,
    8.781799453982851, 1.550013517860879, 1.031249062381747, 1.526929165242378,
    3.422406752555146, 7.964462025926615, 1.150305792701261, 2.766015467833883,
    6.597803992875334, 4.859367503372030,
  -3.216509880131417, 2.906113965081317, 5.862053512785612, 4.468168656522979,
    -1.663731439007003, 2.006191360415653, 6.114556605587009, 5.059283363838881,
    -4.832778328222401, 5.040052435749871, 5.544377368169970, 3.654337461014335,
    6.397673687137877, 3.990761235626036, 1.968069192354027, 4.007185501066716,
    1.590806226463062, -2.041920360224454, 1.972342727051742, 3.371026657168430,
    7.586440734987976, -2.503783744297805, -1.404295330164439, 1.850513531094609,
    3.481356178083440, 3.926524207300429, 5.906618417214159, -3.346656848454868,
    -0.2493135639446889, -1.955296057811105, 8.664457532848232, 1.675496362169158,
    0.8723395253082734, 1.529636995835534, 3.509035347130104, 7.929345249818257,
    1.057667082900209, 2.793155233590146, 6.625375283379160, 5.329178272583427,
  -3.377018169762958, 2.892903119181074, 5.639432825158614, 4.987364755829843,
    -1.441705083849244, 1.977945228432235, 5.647591641274045, 6.105474340188261,
    -4.576921572995084, 5.090057430697018, 4.937760669986710, 3.167176662560316,
    6.323201248117551, 4.102101989782324, 1.190927320502702, 3.893293997714276,
    2.983469908507092, -2.061538334737357, 2.188312658870888, 3.241060230955951,
    7.787024305963874, -2.368717228281943, -1.233328192935760, 1.708010119115257,
    3.098316785398446, 3.782103122907984, 6.035304141205906, -3.295200716566644,
    -0.5643944219683277, -2.223973422041385, 8.647531844513919,
    1.733879868983037, 0.9992853129736721, 1.591389542332374, 3.591316521314882,
    7.881111931339273, 1.037875815410970, 2.887903506806290, 6.653914690103245,
    4.930187556616815,
  -3.243499511813624, 2.861505119635707, 5.547865937084327, 5.054205409391828,
    -1.450026550499627, 2.009569180952303, 5.884022781597032, 5.846291851719477,
    -4.494816816294245, 5.242470795778575, 5.315633915626878, 3.118313930368481,
    6.263501600413233, 4.208433191226665, 1.271889990796535, 3.914066635445268,
    2.827436417263726, -2.067601421779908, 2.247346738924194, 3.437411439824079,
    7.660621823199564, -2.488010855301549, -1.339856783675113, 1.822754170304789,
    3.303919560521436, 3.811683650284884, 6.017681710740752, -3.326905147928402,
    -0.5624001862967027, -2.215401651788850, 8.603763495694775,
    1.740848435821148, 1.098660402379266, 1.669904322937491, 3.650647975603243,
    7.829995673035037, 0.8773861790327103, 2.787337676043454, 6.500316975687538,
    5.409993110220723,
  -3.261101269035726, 2.903872699213573, 5.747234544993702, 4.846248513400098,
    -1.605824048383379, 1.980454974046193, 5.946472146732419, 5.813383580015877,
    -4.543064301680141, 5.266508291927141, 5.287882674267840, 2.930333296282871,
    6.181008835427348, 4.403940393296245, 1.205970402547095, 3.864497681535867,
    2.992906399066627, -2.055379031903006, 2.237072472717980, 3.546159860739998,
    7.662557053630454, -2.600701047713016, -1.215753369411926, 1.773376112913528,
    3.190974555249323, 3.825101636761407, 6.015156737485758, -3.390735214372884,
    -0.1582648304405311, -1.917986863345295, 8.507828594106821, 1.461487971261906,
    0.7995380825702543, 1.600408176257763, 3.702093847396440, 7.979804546288723,
    0.9799853441033393, 2.664757707687734, 6.468143830239463, 5.289411277890451,
  -3.235409117929461, 2.881285947647904, 6.447790177302654, 4.452487852901093,
    -1.893094060216723, 1.524542240146131, 5.752418261017336, 5.999586407200309,
    -3.872279928719233, 5.780136201451364, 5.358493968719256, 2.432023505829708,
    6.289254393699215, 5.546904469729812, 1.502106267059023, 3.633331409711853,
    2.160754860535590, -1.899257293384464, 1.801689556602608, 2.487835779492341,
    8.821849914282101, -1.704609236178317, -1.077258962563566, 2.091787368718893,
    3.291312472791865, 3.960173722753274, 6.086391171891923, -3.444457669313987,
    -0.5114707387184816, -1.758366552048449, 8.718319126081207,
    1.206549723844026, 1.341217333541435, 1.719646361393488, 3.712374669519395,
    7.946937370969962, 1.027871628578638, 2.859292649528902, 6.887503056777743,
    4.785413267041225,
  -3.509820504103284, 2.936120470801730, 5.716925312004083, 5.108481773020319,
    -1.254160946509352, 1.925447637695303, 5.812946483839255, 5.387013942345141,
    -4.863708227886172, 5.031835435840967, 5.039836090427054, 3.041846744036071,
    6.313601220108076, 4.302234071834857, 1.284112482580867, 3.885054925664952,
    2.854933916234350, -2.085655768574008, 2.075314486070811, 2.985015903121788,
    8.010859948487166, -2.194991273525465, -1.232194645060491, 1.671798888738722,
    2.922491798027827, 3.654621348284206, 6.148643695605532, -3.224494799919862,
    -0.7058828277639968, -2.298330104174896, 8.622247943325601, 1.742307082348123,
    1.144446901325226, 1.664378150274813, 3.609316353521339, 7.942899405323680,
    1.141509405849020, 2.781284281048251, 6.529117177837140, 4.694264080813653,
  -3.198583218856307, 2.854978157222592, 5.590713271266168, 4.898686996432050,
    -1.461194527333779, 2.009094449792001, 5.974941123985519, 5.409616955749192,
    -4.806649350791632, 5.071863256299249, 5.305036061670126, 3.247880982317036,
    6.282780635283728, 4.047105690203362, 1.293352478272001, 3.935627965953655,
    2.841802640211119, -2.089947733261740, 2.219337361923091, 3.330172877368538,
    7.739671555794935, -2.400119823193741, -1.356174712494833, 1.799900621559796,
    3.215346686045523, 3.756820411927276, 6.069475746642402, -3.313860296476318,
    -0.5364104462962506, -2.239879779400203, 8.591777810865059, 1.761629851090393,
    1.046857700918966, 1.645471173756973, 3.624742364490974, 7.858003784508190,
    0.9073903660538308, 2.751873742960866, 6.476600022418051, 5.471750722228431 ;

 state_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 state_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 state_postinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 state_postinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 time = 41.666666666666667 ;

 advance_to_time = 41.666666666666667 ;
}
