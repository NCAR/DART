netcdf model_restart {
dimensions:
//	time = UNLIMITED ; 
	t = 5 ;	
	temp = 5 ;
   lat = 180 ;
	lon = 360 ;
variables:
		
	double time(t) ;
	//time:calendar = "none" ;
	//time:units = "days" ;		
	
	double temp(temp) ;
	temp:units = "celsius" ;
   temp:_FillValue = -888888.0 ;
	
	double lat(lat);
	lat:units = "degrees north" ;
   lat:_FillValue = -888888.0 ;
	
	double lon(lon);
	lon:units = "degrees east" ;
   lon:_FillValue = -888888.0 ;
// global attribute
	:title = "garbage lat long for pathological model" ;
	
data:

	time = 0, 1, 2, 3, 4 ;	
	temp = 71.22, 72.314, 73.8872, 10.22, -4.222 ;
	lat = 0, 30, 60, 90, 120 ;
	lon = 0, 60, 120, 180, 240 ;
	//lon = 1, 2, 3 ;	
	//lat = 8, 9, 10 ;
	//lon = 1, 2, 3, 4, 5, 6, 7 ;

}
