netcdf filter_output {
dimensions:
	metadatalength = 64 ;
	member = 40 ;
	time = UNLIMITED ; // (1 currently)
	NMLlinelen = 129 ;
	NMLnlines = 238 ;
	location = 40 ;
variables:
	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "Metadata for each copy/member" ;
	char inputnml(NMLnlines, NMLlinelen) ;
		inputnml:long_name = "input.nml contents" ;
	double time(time) ;
		time:long_name = "time" ;
		time:calendar = "none" ;
		time:units = "days" ;
	double location(location) ;
		location:description = "location coordinates" ;
		location:location_type = "loc1d" ;
		location:long_name = "location on unit circle" ;
		location:storage_order = "X" ;
		location:units = "none" ;
	double state_variable(time, member, location) ;
		state_variable:long_name = "The lorenz-96 wind variables" ;
	double tracer_concentration(time, member, location) ;
		tracer_concentration:long_name = "The lorenz-96 semi lagrangian tracers" ;
	double source(time, member, location) ;
		source:long_name = "The lorenz-96 semi lagrangian tracer sources" ;
	double state_variable_mean(time, location) ;
		state_variable_mean:long_name = "The lorenz-96 wind variables" ;
	double tracer_concentration_mean(time, location) ;
		tracer_concentration_mean:long_name = "The lorenz-96 semi lagrangian tracers" ;
	double source_mean(time, location) ;
		source_mean:long_name = "The lorenz-96 semi lagrangian tracer sources" ;
	double state_variable_sd(time, location) ;
		state_variable_sd:long_name = "The lorenz-96 wind variables" ;
	double tracer_concentration_sd(time, location) ;
		tracer_concentration_sd:long_name = "The lorenz-96 semi lagrangian tracers" ;
	double source_sd(time, location) ;
		source_sd:long_name = "The lorenz-96 semi lagrangian tracer sources" ;
	double state_variable_priorinf_mean(time, location) ;
		state_variable_priorinf_mean:long_name = "The lorenz-96 wind variables" ;
		state_variable_priorinf_mean:units = "unitless" ;
	double tracer_concentration_priorinf_mean(time, location) ;
		tracer_concentration_priorinf_mean:long_name = "The lorenz-96 semi lagrangian tracers" ;
		tracer_concentration_priorinf_mean:units = "unitless" ;
	double source_priorinf_mean(time, location) ;
		source_priorinf_mean:long_name = "The lorenz-96 semi lagrangian tracer sources" ;
		source_priorinf_mean:units = "unitless" ;
	double state_variable_priorinf_sd(time, location) ;
		state_variable_priorinf_sd:long_name = "The lorenz-96 wind variables" ;
		state_variable_priorinf_sd:units = "unitless" ;
	double tracer_concentration_priorinf_sd(time, location) ;
		tracer_concentration_priorinf_sd:long_name = "The lorenz-96 semi lagrangian tracers" ;
		tracer_concentration_priorinf_sd:units = "unitless" ;
	double source_priorinf_sd(time, location) ;
		source_priorinf_sd:long_name = "The lorenz-96 semi lagrangian tracer sources" ;
		source_priorinf_sd:units = "unitless" ;

// global attributes:
		:title = "filter_output.nc" ;
		:assim_model_source = "direct_netcdf_mod.f90" ;
		:creation_date = "YYYY MM DD HH MM SS = 2022 01 06 17 34 07" ;
		:model_source = "$URL$" ;
		:model_revision = "$Revision$" ;
		:model_revdate = "$Date$" ;
		:model = "Lorenz_96_Tracer_Advection" ;
		:model_forcing = 8. ;
		:model_delta_t = 0.05 ;
		:source_rate = 100. ;
		:exponential_sink_folding = 1. ;
		:DART_note = "output prior inflation sd" ;
data:

 MemberMetadata =
  "ensemble member      1                                          ",
  "ensemble member      2                                          ",
  "ensemble member      3                                          ",
  "ensemble member      4                                          ",
  "ensemble member      5                                          ",
  "ensemble member      6                                          ",
  "ensemble member      7                                          ",
  "ensemble member      8                                          ",
  "ensemble member      9                                          ",
  "ensemble member     10                                          ",
  "ensemble member     11                                          ",
  "ensemble member     12                                          ",
  "ensemble member     13                                          ",
  "ensemble member     14                                          ",
  "ensemble member     15                                          ",
  "ensemble member     16                                          ",
  "ensemble member     17                                          ",
  "ensemble member     18                                          ",
  "ensemble member     19                                          ",
  "ensemble member     20                                          ",
  "ensemble member     21                                          ",
  "ensemble member     22                                          ",
  "ensemble member     23                                          ",
  "ensemble member     24                                          ",
  "ensemble member     25                                          ",
  "ensemble member     26                                          ",
  "ensemble member     27                                          ",
  "ensemble member     28                                          ",
  "ensemble member     29                                          ",
  "ensemble member     30                                          ",
  "ensemble member     31                                          ",
  "ensemble member     32                                          ",
  "ensemble member     33                                          ",
  "ensemble member     34                                          ",
  "ensemble member     35                                          ",
  "ensemble member     36                                          ",
  "ensemble member     37                                          ",
  "ensemble member     38                                          ",
  "ensemble member     39                                          ",
  "ensemble member     40                                          " ;

 inputnml =
  "&perfect_model_obs_nml                                                                                                           ",
  "   read_input_state_from_file = .false.,                                                                                         ",
  "   single_file_in             = .true.                                                                                           ",
  "   input_state_files          = \"perfect_input.nc\"                                                                               ",
  "                                                                                                                                 ",
  "   write_output_state_to_file = .true.,                                                                                          ",
  "   single_file_out            = .true.                                                                                           ",
  "   output_state_files         = \"perfect_output.nc\"                                                                              ",
  "   output_interval            = 1,                                                                                               ",
  "                                                                                                                                 ",
  "   async                      = 0,                                                                                               ",
  "   adv_ens_command            = \"./advance_model.csh\",                                                                           ",
  "                                                                                                                                 ",
  "   obs_seq_in_file_name       = \"obs_seq.in\",                                                                                    ",
  "   obs_seq_out_file_name      = \"obs_seq.out\",                                                                                   ",
  "   init_time_days             = 0,                                                                                               ",
  "   init_time_seconds          = 0,                                                                                               ",
  "   first_obs_days             = -1,                                                                                              ",
  "   first_obs_seconds          = -1,                                                                                              ",
  "   last_obs_days              = -1,                                                                                              ",
  "   last_obs_seconds           = -1,                                                                                              ",
  "                                                                                                                                 ",
  "   trace_execution            = .false.,                                                                                         ",
  "   output_timestamps          = .false.,                                                                                         ",
  "   print_every_nth_obs        = -1,                                                                                              ",
  "   output_forward_op_errors   = .false.,                                                                                         ",
  "   silence                    = .false.,                                                                                         ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&filter_nml                                                                                                                      ",
  "   single_file_in               = .true.,                                                                                        ",
  "   input_state_files            = \'filter_input.nc\'                                                                              ",
  "   input_state_file_list        = \'\'                                                                                             ",
  "                                                                                                                                 ",
  "   stages_to_write  = \'preassim\', \'analysis\', \'output\'                                                                           ",
  "                                                                                                                                 ",
  "   single_file_out              = .true.,                                                                                        ",
  "   output_state_files           = \'filter_output.nc\'                                                                             ",
  "   output_state_file_list       = \'\'                                                                                             ",
  "                                                                                                                                 ",
  "   output_interval              = 1,                                                                                             ",
  "   output_members               = .true.                                                                                         ",
  "   num_output_state_members     = 20,                                                                                            ",
  "   output_mean                  = .true.                                                                                         ",
  "   output_sd                    = .true.                                                                                         ",
  "                                                                                                                                 ",
  "   ens_size                     = 40,                                                                                            ",
  "   num_groups                   = 1,                                                                                             ",
  "   perturb_from_single_instance = .true.,                                                                                        ",
  "   perturbation_amplitude       = 0.2,                                                                                           ",
  "   distributed_state            = .true.                                                                                         ",
  "                                                                                                                                 ",
  "   async                        = 0,                                                                                             ",
  "   adv_ens_command              = \"./advance_model.csh\",                                                                         ",
  "                                                                                                                                 ",
  "   obs_sequence_in_name         = \"obs_seq.out\",                                                                                 ",
  "   obs_sequence_out_name        = \"obs_seq.final\",                                                                               ",
  "   num_output_obs_members       = 20,                                                                                            ",
  "   init_time_days               = 0,                                                                                             ",
  "   init_time_seconds            = 0,                                                                                             ",
  "   first_obs_days               = -1,                                                                                            ",
  "   first_obs_seconds            = -1,                                                                                            ",
  "   last_obs_days                = -1,                                                                                            ",
  "   last_obs_seconds             = -1,                                                                                            ",
  "                                                                                                                                 ",
  "   inf_flavor                  = 2,                       0,                                                                     ",
  "   inf_initial_from_restart    = .false.,                 .false.,                                                               ",
  "   inf_sd_initial_from_restart = .false.,                 .false.,                                                               ",
  "   inf_deterministic           = .true.,                  .true.,                                                                ",
  "   inf_initial                 = 1.0,                     1.0,                                                                   ",
  "   inf_lower_bound             = 1.0,                     1.0,                                                                   ",
  "   inf_upper_bound             = 1.2,                     1.2,                                                                   ",
  "   inf_damping                 = 0.9,                     1.0,                                                                   ",
  "   inf_sd_initial              = 0.6,                     0.0,                                                                   ",
  "   inf_sd_lower_bound          = 0.6,                     0.0,                                                                   ",
  "   inf_sd_max_change           = 1.05,                    1.05,                                                                  ",
  "                                                                                                                                 ",
  "   trace_execution              = .false.,                                                                                       ",
  "   output_timestamps            = .false.,                                                                                       ",
  "   output_forward_op_errors     = .false.,                                                                                       ",
  "   write_obs_every_cycle        = .false.,                                                                                       ",
  "   silence                      = .false.,                                                                                       ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&smoother_nml                                                                                                                    ",
  "   num_lags              = 0,                                                                                                    ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .false.,                                                                                              ",
  "   restart_in_file_name  = \'smoother_ics\',                                                                                       ",
  "   restart_out_file_name = \'smoother_restart\'                                                                                    ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&ensemble_manager_nml                                                                                                            ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&assim_tools_nml                                                                                                                 ",
  "   filter_kind                     = 1,                                                                                          ",
  "   cutoff                          = 0.2,                                                                                        ",
  "   sort_obs_inc                    = .false.,                                                                                    ",
  "   spread_restoration              = .false.,                                                                                    ",
  "   sampling_error_correction       = .false.,                                                                                    ",
  "   adaptive_localization_threshold = -1,                                                                                         ",
  "   output_localization_diagnostics = .false.,                                                                                    ",
  "   localization_diagnostics_file   = \'localization_diagnostics\',                                                                 ",
  "   print_every_nth_obs             = 0,                                                                                          ",
  "   rectangular_quadrature          = .true.,                                                                                     ",
  "   gaussian_likelihood_tails       = .false.,                                                                                    ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&cov_cutoff_nml                                                                                                                  ",
  "   select_localization = 1,                                                                                                      ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&reg_factor_nml                                                                                                                  ",
  "   select_regression    = 1,                                                                                                     ",
  "   input_reg_file       = \"time_mean_reg\",                                                                                       ",
  "   save_reg_diagnostics = .false.,                                                                                               ",
  "   reg_diagnostics_file = \"reg_diagnostics\",                                                                                     ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&obs_sequence_nml                                                                                                                ",
  "   write_binary_obs_sequence = .false.,                                                                                          ",
  "   read_binary_file_format   = \'native\'                                                                                          ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&obs_kind_nml                                                                                                                    ",
  "   assimilate_these_obs_types = \'\'# \'RAW_STATE_VARIABLE\',                                                                        ",
  "\t\t\t\t#\'RAW_TRACER_CONCENTRATION\',                                                                                                 ",
  "\t\t\t\t#\'RAW_TRACER_SOURCE\'                                                                                                         ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&model_nml                                                                                                                       ",
  "   model_size        = 120,                                                                                                      ",
  "   forcing           = 8.00,                                                                                                     ",
  "   delta_t           = 0.05,                                                                                                     ",
  "   time_step_days    = 0,                                                                                                        ",
  "   time_step_seconds = 3600,                                                                                                     ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&utilities_nml                                                                                                                   ",
  "   termlevel      = 1,                                                                                                           ",
  "   module_details = .false.,                                                                                                     ",
  "   logfilename    = \'dart_log.out\',                                                                                              ",
  "   nmlfilename    = \'dart_log.nml\',                                                                                              ",
  "   write_nml      = \'file\',                                                                                                      ",
  "   print_debug    = .false.,                                                                                                     ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&mpi_utilities_nml                                                                                                               ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&preprocess_nml                                                                                                                  ",
  "   overwrite_output        = .true.                                                                                              ",
  "   input_obs_def_mod_file  = \'../../../observations/forward_operators/DEFAULT_obs_def_mod.F90\'                                   ",
  "   output_obs_def_mod_file = \'../../../observations/forward_operators/obs_def_mod.f90\'                                           ",
  "   input_obs_qty_mod_file  = \'../../../assimilation_code/modules/observations/DEFAULT_obs_kind_mod.F90\'                          ",
  "   output_obs_qty_mod_file = \'../../../assimilation_code/modules/observations/obs_kind_mod.f90\'                                  ",
  "   obs_type_files          = \'../../../observations/forward_operators/obs_def_1d_state_mod.f90\'                                  ",
  "   quantity_files          = \'../../../assimilation_code/modules/observations/oned_quantities_mod.f90\'                           ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&obs_sequence_tool_nml                                                                                                           ",
  "   filename_seq      = \'obs1.out\', \'obs2.out\',                                                                                   ",
  "   filename_seq_list = \'\',                                                                                                       ",
  "   filename_out      = \'obs_seq.combined\',                                                                                       ",
  "   first_obs_days    = -1,                                                                                                       ",
  "   first_obs_seconds = -1,                                                                                                       ",
  "   last_obs_days     = -1,                                                                                                       ",
  "   last_obs_seconds  = -1,                                                                                                       ",
  "   print_only        = .false.,                                                                                                  ",
  "   gregorian_cal     = .false.,                                                                                                  ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&obs_diag_nml                                                                                                                    ",
  "   obs_sequence_name     = \'obs_seq.final\',                                                                                      ",
  "   bin_width_days        = -1,                                                                                                   ",
  "   bin_width_seconds     = -1,                                                                                                   ",
  "   init_skip_days        = 0,                                                                                                    ",
  "   init_skip_seconds     = 0,                                                                                                    ",
  "   Nregions              = 3,                                                                                                    ",
  "   trusted_obs           = \'null\',                                                                                               ",
  "   lonlim1               = 0.00, 0.00, 0.50                                                                                      ",
  "   lonlim2               = 1.01, 0.50, 1.01                                                                                      ",
  "   reg_names             = \'whole\', \'lower\', \'upper\'                                                                             ",
  "   create_rank_histogram = .true.,                                                                                               ",
  "   outliers_in_histogram = .true.,                                                                                               ",
  "   use_zero_error_obs    = .false.,                                                                                              ",
  "   verbose               = .false.                                                                                               ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&schedule_nml                                                                                                                    ",
  "   calendar        = \'Gregorian\',                                                                                                ",
  "   first_bin_start =  1601,  1,  1,  0,  0,  0,                                                                                  ",
  "   first_bin_end   =  2999,  1,  1,  0,  0,  0,                                                                                  ",
  "   last_bin_end    =  2999,  1,  1,  0,  0,  0,                                                                                  ",
  "   bin_interval_days    = 1000000,                                                                                               ",
  "   bin_interval_seconds = 0,                                                                                                     ",
  "   max_num_bins         = 1000,                                                                                                  ",
  "   print_table          = .true.                                                                                                 ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&obs_seq_to_netcdf_nml                                                                                                           ",
  "   obs_sequence_name = \'obs_seq.final\',                                                                                          ",
  "   obs_sequence_list = \'\',                                                                                                       ",
  "   append_to_netcdf  = .false.,                                                                                                  ",
  "   lonlim1    =    0.0,                                                                                                          ",
  "   lonlim2    =    1.0,                                                                                                          ",
  "   verbose    = .true.                                                                                                           ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&state_vector_io_nml                                                                                                             ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&quality_control_nml                                                                                                             ",
  "   input_qc_threshold       =  3.0,                                                                                              ",
  "   outlier_threshold        = -1.0,                                                                                              ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&integrate_model_nml                                                                                                             ",
  "   trace_execution = .true.                                                                                                      ",
  "   ic_file_name    = \'temp_ic.nc\'                                                                                                ",
  "   ud_file_name    = \'temp_uc.nc\'                                                                                                ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "&model_mod_check_nml                                                                                                             ",
  "  input_state_files     = \'perfect_input.nc\'                                                                                     ",
  "  output_state_files    = \'mmc_output.nc\'                                                                                        ",
  "  num_ens               = 1                                                                                                      ",
  "  single_file           = .false.                                                                                                ",
  "  test1thru             = 0                                                                                                      ",
  "  run_tests             = 1,2,3,4,5,6,7                                                                                          ",
  "  x_ind                 = 2                                                                                                      ",
  "  loc_of_interest       = 0.3                                                                                                    ",
  "  quantity_of_interest  = \'QTY_STATE_VARIABLE\'                                                                                   ",
  "  interp_test_dx        = 0.02                                                                                                   ",
  "  interp_test_xrange    = 0.0, 1.0                                                                                               ",
  "  verbose               = .true.                                                                                                 ",
  "  /                                                                                                                              " ;

 time = 49.9583333333333 ;

 location = 0, 0.025, 0.05, 0.075, 0.1, 0.125, 0.15, 0.175, 0.2, 0.225, 0.25, 
    0.275, 0.3, 0.325, 0.35, 0.375, 0.4, 0.425, 0.45, 0.475, 0.5, 0.525, 
    0.55, 0.575, 0.6, 0.625, 0.65, 0.675, 0.7, 0.725, 0.75, 0.775, 0.8, 
    0.825, 0.85, 0.875, 0.9, 0.925, 0.95, 0.975 ;

 state_variable =
  1.82825739350251, 7.5938903016588, 5.04840911731483, -5.17914273362721, 
    1.46884352186564, 4.11570872948408, 8.47408470831022, 4.15017459318918, 
    -1.59597992633523, -0.519290585451951, 0.410641152695634, 
    2.58968782642916, 6.86073421733203, 1.06033564575766, 3.19325037121091, 
    4.44190719411893, 6.06828145816484, -1.80190723107405, 
    -0.0820399554152673, -1.74844552242657, 7.47727356044064, 
    3.22535441173144, -1.54447809301826, 0.440102854408848, 8.90218809094372, 
    3.24927114737404, -1.36117119695556, 0.471694625532235, 
    0.432336235465306, 5.11364590054238, 4.14471082071672, -2.43576214643811, 
    1.90560185730282, 11.2107783029596, -0.0801984609855013, 
    3.11899881106735, 5.55306251235197, 4.57840459968543, -1.11362562629826, 
    -1.04314024556569,
  5.52526804329785, 3.61481037192371, 3.97993195464659, 0.556802440330242, 
    -3.94191810500834, 2.47888464849376, 4.32818625737223, 6.19424410329768, 
    -0.705223681032597, -3.22323440260423, 1.25580022829852, 
    3.35994946562654, 9.81544831151799, 7.06820817380818, 0.959122181865746, 
    3.9967377646026, -1.90028305053486, -0.597306784997154, 
    0.606484079432262, 7.53992951253058, -1.2441697227289, -5.52077884222918, 
    1.28769425837758, 1.84195273074883, 8.41125893872542, 4.09315586733171, 
    -2.47854936959215, 2.90255624988894, 2.56405704600802, 5.0240952116887, 
    8.46922260081886, -1.92091016779032, 2.2746687814619, 1.75903107532989, 
    0.0584708024013069, 0.801315435303813, 7.27596079351922, 
    -0.653418069368405, -2.9940548276682, 2.40720296237393,
  5.06239052187456, 4.43432813258343, 7.47955710523757, 5.06274898435458, 
    -2.09657350644547, 1.68421490567551, 2.54392749592549, 0.794462655262644, 
    3.06361316977842, 10.0776442454613, 1.37640763258809, 0.0814905131038705, 
    3.93199635410117, 2.07463373562359, 4.11908878477941, 6.62327684935105, 
    0.688689804970698, -4.19027840623471, 1.63783409351106, 3.89251218535814, 
    7.75164977353037, 1.78167987287189, -3.65201088086235, 0.606691107390003, 
    5.57081813345366, 8.34902450197484, -0.724173647707681, 
    0.122462456869957, -1.26022101507113, 1.10954394812522, 5.62514315528083, 
    11.4103892898948, 3.70984788311416, 2.6960092534059, 6.87184235873404, 
    -1.44820711120444, -3.94956366709169, -0.7200215723552, 
    -1.86211493981668, 3.5523089202296,
  0.902025561832744, -1.64162903154639, -3.11962063651157, 
    -0.994160246284155, -3.37436046856884, 2.43005801739715, 
    8.75614173344054, -1.71602551981352, 2.23846670698898, 6.49673557241401, 
    2.34917105479758, -0.257184044692599, 4.06340097597292, 9.43393438260215, 
    -1.89710770648213, 1.81796520270031, 0.606910761483172, 
    -0.236870081495473, 1.09632962945094, 4.7725772322631, 6.09927415917005, 
    -2.20846871292985, -1.98866898902934, -0.824053240860295, 
    0.673402594205652, 7.73127964522868, 4.27258486070095, -4.82781539131029, 
    1.29957677494494, 6.48758905044165, 4.90750828877434, 
    -0.0670568300412724, 5.50030113312845, 9.78631480100078, 
    4.12742480939089, 4.15795804726526, 1.92624618290053, -1.0658445103156, 
    3.71673432756463, 8.82922778198363,
  8.89102423470524, -1.7770663124641, 3.0637867084599, 2.5661231038593, 
    5.07118799096199, 7.87081766727141, -1.22293862218312, -1.34438953216367, 
    -1.00480998716153, 0.684757404163928, 3.44700868068801, 7.00118446116095, 
    0.0261513251382459, 2.21350080888596, 6.93224390161412, 7.86492387396317, 
    -0.764450407146411, 3.88417802455718, 8.7750932637475, 4.81616836942899, 
    -0.946763313938641, 0.347391794761807, 5.90905314420361, 
    8.06123448564217, -4.68954080465979, 2.93131132273522, 1.70642301284029, 
    6.07030936009015, 0.983919404736096, -1.92996437578317, 2.0511359168855, 
    10.0826431844775, 6.28669909756843, 3.56506030856137, 4.27875404234006, 
    1.06109216109558, 3.70489569152756, 2.18176229967264, 0.775513618786849, 
    3.91554502292307,
  -3.59037481326941, -0.103551540778414, 9.67066736114967, 1.0329641788617, 
    -1.54018566072783, -1.2565657985965, 3.06361367408572, 5.92126693749055, 
    4.57878337862373, -3.48368672228484, -1.67483366635272, 
    -2.70009386658155, 5.4385174171984, 6.70965936755244, 1.59468213072878, 
    4.61136169838767, 8.04077562343543, 0.079788225617146, 
    -0.165525889821838, 5.38270291756546, 5.06186753513287, 
    -2.91321390901998, 4.19588159566729, 4.9231796274774, 2.63611166127997, 
    4.56390508906448, 5.13855727751081, -0.259588892447064, 3.41505115861375, 
    5.90394393449218, 0.87878148618223, -3.5941787251606, 1.79643821279539, 
    2.63691353292546, 6.62377109259681, 2.09895172495233, -4.1822001855837, 
    0.938254924730014, 5.22612650448232, 0.994091849022955,
  2.71745911588437, 5.81812608268125, 8.47840734760387, 0.782950617095143, 
    2.49727291878279, 1.54458326915192, 2.68408002774065, 6.88313419010329, 
    1.12064707825847, -5.32230329793631, 4.03345828469534, 3.62220514378907, 
    2.6679712434918, 7.1717398282501, 5.96034060523945, 3.70534409651877, 
    4.77398292868482, -0.609041745121553, -1.06642203106336, 
    0.875268040710253, 6.29335844586117, 1.86267748001819, -1.77771771677295, 
    4.04562188036428, 7.71518592695659, 2.85186570035023, 2.93934295230837, 
    -0.719875012542152, -0.969877937422995, 0.246673068250398, 
    7.68962121072684, -0.543383567646832, -3.18247120308426, 
    0.594292052747149, 1.94627361755255, 6.26735836635197, -1.27963378822067, 
    -3.8499123460927, 2.38039570663181, 3.83835376269132,
  2.50344279896712, 8.66423449508454, 7.57093033656499, 1.71967075399183, 
    2.23237378025595, 2.66074129957041, -2.02383878461068, 
    0.0448537816071762, 0.300238855062496, 4.7133107160052, 9.49716330280643, 
    2.33587998733134, 3.57027667952259, 3.59138929101437, -3.3054473818952, 
    2.57218517267577, 10.005248056995, -1.30170910935642, 0.241220277919142, 
    3.44705931377125, 10.4307730953837, -0.635129628271661, 1.05858042022168, 
    3.09077174574447, -0.175703724079194, 3.26248797350594, 7.74515940874136, 
    4.20761966751902, -2.47878850969681, -1.34800454536332, 3.16652614678792, 
    8.94976229807271, 3.13633876533214, -1.49515044056822, -4.55626494153391, 
    2.39879385352423, 4.97050566743283, 4.34988722085772, 2.4851421020715, 
    -2.74873960963628,
  0.0447778766464132, -0.598147925709112, 2.18798247737252, 5.76278101669324, 
    0.898754095938541, 2.05140554034146, 4.14403194085018, 2.47877459549506, 
    3.3233066667325, 7.76390202582411, -1.66836661838544, 2.4998971666213, 
    2.06565045315491, 6.2008011681781, 4.70718744274896, -4.11363938626985, 
    4.76706740460298, 1.98832814927344, 1.55854489560045, 0.336471205996539, 
    4.91460265040302, 3.13488664605301, -3.32943280990085, 0.253871312140409, 
    4.90924974559555, 6.3140127371184, -0.143928547040003, 4.20761083920496, 
    6.29428887242308, -2.94735136612336, 1.80870244851633, 6.29360835270399, 
    6.14153657391907, -3.99195533347243, 7.0327423915333, 0.518400107943933, 
    -0.404204981088641, 3.8186578744554, 10.4102716399596, -3.10266439577525,
  5.08216711217846, 10.3236074820639, -0.236065644532693, -0.907797951233902, 
    4.37827667340295, 0.155230917252598, 1.03754952410846, 1.24669357171698, 
    3.33805763795605, 6.23341280058172, 3.55556867266729, -3.16052508292429, 
    -2.91048873379752, 1.08952764006476, 4.42817198786124, 6.20640744344399, 
    -0.199758946864091, -0.785505174801257, 1.70793943641414, 
    10.1221294473987, 5.87505301221021, 3.72270583527055, 7.3200192796136, 
    2.71386292579198, -2.02344851054871, -1.9836840839321, 
    -0.421163355989692, 8.49623613755782, 1.56241037591188, 
    0.422570625349998, 5.6025534883531, 8.15301959306537, -1.37190392566508, 
    5.40803394792671, 3.72422368923785, 1.45547506646353, 2.71883034308865, 
    6.4366273818399, 3.12232393620469, 1.27715791730602,
  -1.16736982712279, 10.5368286300181, 2.39378232309306, -2.77441702189993, 
    0.732735476421828, 5.65980122749321, 4.28839529844636, -1.37675800746328, 
    2.64195502698183, 10.0897572227836, -3.95378453694914, 1.78404839806502, 
    1.94067782715895, 10.1289812501007, 0.820481329865637, -3.59739687228466, 
    1.23897280990939, 3.45071126665519, 5.43735948288978, -0.819137654243359, 
    0.412049418637937, 1.22088999900356, 7.49519344895353, 1.35912668057932, 
    2.35037086834509, 4.92817637270889, 5.82793088327345, -2.25941609706977, 
    -2.86893304331117, -1.058543874956, 0.700818277859562, 3.12283116749832, 
    7.34149085607751, -1.15531598587724, 2.12231481832949, 2.66477041839764, 
    4.02758566900611, 6.50439562152082, -3.53620745516544, -1.81611132966477,
  -1.12308810177214, 3.48033524891586, 5.27976111279035, -5.35052089868444, 
    0.845904552189998, 0.502768835645749, 5.89244517732684, 3.40728863903612, 
    -2.85072292197416, 2.02568942572951, 1.58939966302106, 6.56981798363781, 
    1.00567123098804, 0.636790733844825, 1.30614743543499, 5.49060231488577, 
    0.835553835115192, -3.55217558698586, 2.33476353877811, 8.30977529710938, 
    5.37373445897983, -2.51204749706263, 0.898241041548106, 1.8018024954296, 
    9.03379501651533, 0.432017378182092, -2.77485760691741, 2.14768911426091, 
    9.21200499613669, -0.968370663174193, 0.444214775663629, 
    1.99829499216996, 6.90144332945681, 0.189211701331351, -2.79209576178731, 
    4.16434817568388, 4.17832674814001, 1.5656291438309, 6.92126294897802, 
    3.64828524429692,
  9.64342690455948, 1.54714668108153, 4.98859466639001, 3.69446471049993, 
    3.11066964211861, 3.11850598122865, -2.37624418233903, 1.49621213980459, 
    2.29912854177667, 6.48197040351819, -2.61381217389488, -3.11173094910203, 
    -0.599822733494239, 2.5597012308796, 6.33313348190561, 1.32426513665419, 
    3.1427792477199, 7.77928428443633, 1.03353759934569, -4.00562789472345, 
    2.43434630780361, 9.8275227948172, 3.73865809577877, 1.61001881962201, 
    1.23872324072645, -2.192101090003, 1.48115347537371, 4.48908995648253, 
    7.93993803613821, 2.3880051845137, 4.08934777844313, 7.97349959772967, 
    5.86259271309261, 2.50680513601125, 1.13020007592294, 1.56464868118252, 
    5.91411426434443, 3.19025546739495, -0.827462165664302, 6.84128812230109,
  6.20021010904294, 5.2737282054692, -6.65674348348413, 2.28382619593925, 
    3.16559652902957, 5.38459847711465, -0.688373197428854, 1.45703367030741, 
    2.88711793688753, 8.33363974669149, -3.67348467398405, 
    -0.588720964512214, -1.74445781442207, 7.3726735333734, 
    -1.09885892092734, -0.730773298763309, -1.31434488106449, 
    8.03308217253148, -0.518107374199921, -2.59242114226947, 
    0.710126431066017, 3.6731096232335, 9.27994539658595, -5.24044316222712, 
    1.44898397729805, 1.97018326027656, 5.60309945298253, 0.0891412862004906, 
    1.8858631197993, 6.36639109871364, 8.1296663932737, -2.11286493780026, 
    1.96992371896987, 3.18903766170516, 0.615493029856567, 2.67618320508996, 
    6.12014734799494, -2.19511717150999, -1.91481966690138, -0.093334443265763,
  1.78421135128605, 7.80736325873595, -2.29201239994014, -2.05812709726036, 
    0.691352364293608, 3.31536421950906, 6.16555301929759, 4.34689506879737, 
    -2.47732733205512, -0.110491007427653, 3.69752264412479, 
    8.36721625931876, -0.139319494266469, 1.00458972814011, 
    -1.14155834018265, 1.87528482719122, 4.66182899767224, 8.08770688681352, 
    0.430142768259464, -2.51632303591917, 2.60538611696439, 7.80820189848057, 
    -1.16439032995587, -0.147802659566093, 2.53673261951989, 
    9.94520431456408, -2.44317745668789, -1.70438307685708, 
    0.292926666952215, 7.69502910580835, 5.67952823604219, 1.75775414252878, 
    3.85475143516498, 1.42450766682757, -1.24633186928836, 1.52326436045509, 
    -1.60742127309982, 3.52548405017137, 4.85238222022089, -3.6365583860058,
  1.76104647804631, 2.19545910038938, 4.76579636395886, 8.16472454997188, 
    -4.1498377396874, 1.46466193247344, 4.78153133745566, 5.14397149882012, 
    4.30071804116359, 5.60880534834948, -0.313653016391514, 
    -4.62418572848228, 1.24941787217604, 3.62244892234034, 11.2343888692272, 
    0.0839962985077481, 0.677043932233121, 2.53291412274605, 
    1.35977758484124, 2.5266713289795, 9.92729134261537, 4.15323013084148, 
    0.753036303018856, 0.531599068210203, 3.19125407750626, 6.92746703982962, 
    1.80251967876913, 3.28688231144162, 7.68375957090126, 1.66670091771936, 
    -2.3159407971991, 2.88447783279423, 7.60863653198746, -2.71073740422608, 
    -1.05344427988629, -1.11594337652951, 0.763993478713327, 
    3.21114264996626, 8.54462587650543, -0.458375071094483,
  3.60933454822814, 4.26597796812268, -1.36033115263818, 2.18552832271237, 
    4.53278038742335, 10.1876663062858, 4.60879757858018, -5.08123533346925, 
    4.09192757265664, 8.38112819897418, -2.38005290434575, 2.05363481427547, 
    4.46977418081237, 4.80784380877924, 1.42723780640545, 4.1358897569151, 
    8.09177519300417, -1.04061843469118, -4.8487738547827, -1.19096372886621, 
    4.20860706459932, 5.75732215711915, 2.04389314570499, 4.17475525691036, 
    5.58719543799104, -0.174353392758563, -0.907821713760702, 
    3.7712599822451, 10.7684190619661, 6.71083817022442, 0.679775593486533, 
    0.539533109604533, 4.06877841290198, 2.50525104624228, 1.04966796526419, 
    4.12017122248525, 7.95536226052906, 3.4967818780758, 5.38585513719996, 
    5.98803113373873,
  3.37339822915794, -1.62954560106241, -1.46762366382958, 7.77475050012251, 
    6.23782732463135, -2.8447442940634, 1.90946648020335, 2.16494216220442, 
    4.03040806048984, 3.78356969064354, -2.56333284589955, 3.16950687227215, 
    6.22971981078778, 5.84084783328358, 6.29369233464385, 2.02963634521039, 
    -0.55052674365415, 4.66607241057798, 10.1814675135431, -1.74520682205487, 
    0.0550977126976827, -0.0135333898661182, 0.711843950800448, 
    3.4411427686808, 10.3618458933292, 0.642888945787452, 1.96741989107809, 
    5.28302267203385, -0.299787434870699, 3.76055098293409, 4.35635321655087, 
    6.25934046743885, -2.68293480896093, -0.927364341741067, 
    -0.374678376240016, 2.50198920506727, 8.50053268580746, 
    -1.88803487390582, 0.0254344137302127, -1.93112229994697,
  -2.27047806856358, 2.02531530938923, 7.38351453062748, 6.84781309679847, 
    3.72628551007967, -0.270405505951246, 3.73096066907231, 4.29849892498318, 
    4.65752434845729, 4.91623214371043, -3.36700533987486, 
    -0.182834446064756, 0.37035362602329, 2.74828466571555, 7.57229019142634, 
    -1.5308763679946, -5.24246714244677, -1.48452729974483, 6.81681597777433, 
    3.61161510484049, 1.22381933600875, 5.44964122693215, 7.28716329172089, 
    1.79074434080345, 4.03686405734802, 2.23719396847641, -4.50632971412232, 
    4.61181720496056, 6.30635246361062, 4.13530716366867, 3.66313136591096, 
    -0.113276557989663, 5.98123116882995, 3.07696538709957, 
    0.365866219901421, 4.50562653576722, 10.8023420254096, 0.582475042359806, 
    1.46137265332981, 0.822104642214174,
  -1.16071028493993, -1.08015344998413, 4.34543616328896, 3.366857846623, 
    1.26108456494128, 2.2073857199258, 4.38247896576575, 5.14950468719358, 
    -6.07608898341324, 4.93929752919902, -2.2275217154032, 4.98997557625196, 
    4.9877358335437, -7.09096265823603, 3.41354238723238, 5.77515420510488, 
    4.58304049627976, 4.85571348548236, 0.0617333399669033, 
    -4.82723487172037, 1.99405923368094, 1.23617318139615, 4.59134179935578, 
    9.2293593473917, 2.07572037837234, -0.529575630485357, -0.90011827473682, 
    0.158213434965956, 5.30145328767026, 8.48941996103061, 
    -0.694065553118269, 3.55800917819427, 0.348929650362396, 
    0.424981505936087, 1.70147768837023, 9.21937062526089, 1.92666686411184, 
    -3.02453062983829, 2.02976085049252, 9.45212674256847,
  -0.130990995498365, -3.92124999725735, 1.02289666421947, 7.71363396049351, 
    5.73244280220291, 0.378107670532572, -1.49209556076639, 
    -3.37865599373499, 1.79860945402345, 2.7933924024144, 5.75454392986089, 
    7.40215722521069, 2.01929205405562, 4.5277183320539, 2.55416646723952, 
    -4.38347685099994, 1.21182832048626, 7.80389528728718, 6.23483681683618, 
    -1.53885975955847, 5.26439575965929, 5.2923804908074, 1.36976754369074, 
    3.33854658496024, 5.405869116365, 1.41145852134172, -2.69894129598122, 
    0.96620917770655, 2.71430519442524, 7.91464776313223, -2.38643117430021, 
    -1.38177885996912, -0.382155554605311, 4.39321314122949, 
    8.60418088911479, 1.42662994327554, 4.8676489453119, 4.38414064253163, 
    3.19276505520845, 4.94510481435672,
  1.82228839625586, 9.05453591138202, -1.14882453949824, 1.11132624497894, 
    -0.688300647330676, 1.059841156173, 0.900367907651795, 1.73111322904073, 
    5.24335889941847, 4.15606424133042, -4.81119425133298, 1.29077441640566, 
    2.74452169065188, 8.68225709457463, 4.35498728684485, -1.82759632040219, 
    0.457271665907449, 0.443748804688058, 3.33805862074967, 6.73352877646884, 
    -3.51341934538032, 2.94908733416597, 1.54579078489833, 1.02616180543571, 
    6.15541551881646, 12.5535186158069, -0.140128468046894, 3.47850510428026, 
    3.73573493783793, -0.453565714684684, 4.12446016127282, 7.84954335651151, 
    7.50790132772668, 5.28918144479095, 0.568977996556383, 3.74688144182495, 
    7.0601305076602, -1.52187567797238, -2.0093273662355, -0.556892935068328,
  2.73477456369622, 3.81836132944473, 4.62350239191216, -4.04886209483087, 
    -0.0781357101766978, 2.70090339591741, 5.83745297987014, 
    3.72940596382458, 3.60514380144625, -3.00366890402372, 
    -0.449354110500914, -2.96558478644174, 5.34003272133493, 
    2.19204545637979, -2.50810640863344, 3.26473693535143, 7.95701927145493, 
    5.23345041352083, 7.04540056560078, 5.83777756029058, 0.308455900479413, 
    5.14365739092805, 8.2951317126684, 4.16690726423259, 2.01042941869113, 
    -1.58562899095266, -0.794026156425409, 4.62381488281325, 
    4.71002362343893, -0.0810872397500647, 3.03556106521619, 
    6.91540639589406, -3.5904915377252, 1.46700663382709, 1.88515458412311, 
    2.8909680694277, 4.09698583993485, 3.69321953062362, -4.91991239929011, 
    3.93372408134448,
  0.898416372268932, 4.00390243936033, 8.19442728254305, 1.78863230950993, 
    -6.92021374686626, 0.0761834065157725, -1.61094235513106, 
    3.4576607348263, 7.72568670149097, -2.40003602021453, 4.39749080189046, 
    6.99840298127122, 4.3193340797823, 1.64141084643696, 3.26635780815097, 
    5.10161080256063, -1.32705094652356, -3.47498675157133, 2.2020155305458, 
    6.40607016112471, 4.10151273180017, -0.851199641809621, 
    -2.58521889778043, 0.643916966626015, 11.5474600407099, 4.76639314889466, 
    -0.968225764766969, 0.83858941034999, 1.9676105547231, 6.57429834479061, 
    4.50453059212582, 0.670011916306604, 5.09140211673065, 5.40291979457795, 
    -0.617654806530146, 4.86412186919177, 8.38916153013165, 2.15163580258782, 
    -0.402617400335147, -3.66560428604886,
  1.80891472192322, 7.00481346739432, 7.52523943194725, 2.68327334970647, 
    2.59759271610131, -5.14057893271644, -0.275171649442602, 
    -2.46140322051566, 2.48787428245215, 10.2205683843669, 0.505800311934223, 
    3.0571204746988, 5.11829075126808, -1.9299039679581, 0.892159290589246, 
    -0.871326706234923, 6.74784019879947, 3.76653441555623, 
    -2.08540530621182, 2.25664080107708, 6.35659039746194, 
    -0.607399359594481, 2.18808924352984, 7.01389669366115, 
    -0.0971779450300117, 1.84751507610505, 0.8161696563461, 6.95672848674862, 
    -2.32654949649563, -1.37527302679012, -5.72039697632681, 
    2.17812564229488, 2.38035326609107, -4.6607472407563, 1.28729305620323, 
    6.27748008531271, 4.37952520291574, 1.62809678334821, -4.92080543200426, 
    2.46132838872904,
  6.51548676489146, 4.53326061881859, -3.87942441806006, -2.18559609647723, 
    -0.0609028200577152, 9.09144414223821, 3.55542234395244, 
    -1.78002023258517, -0.350667993542292, -0.321120150381812, 
    -0.159279769535703, 7.17156885940749, 2.07982291539714, -1.4055168911577, 
    3.93418247010863, 10.6550601608433, 6.61799436846947, 5.11503738971413, 
    4.39481595888422, 2.92676011699812, 7.62272206725922, 7.58926566456918, 
    0.515778187478299, 4.7973360360155, 5.28842518118127, 2.13498127906221, 
    4.67884867423293, 0.293145688959895, -0.50464837333353, 0.97430922351386, 
    8.63822996894834, -0.620346339557031, 3.45877924698455, 
    0.288519020664128, 0.658414978482274, 9.89491043792493, 2.02731013025125, 
    -2.23618072579149, 1.93600851827565, 4.44543726522893,
  -3.59983479266975, 3.71697169532688, 5.00192747352454, 1.88631465399381, 
    5.91700932227147, 5.41403165656923, -2.97927970967409, 3.03750504892774, 
    7.13650078572688, 2.91666981554828, -3.47735217787243, 0.164932352146481, 
    1.83474530976769, 7.31470981644416, -0.228246064547092, 3.10977425843199, 
    8.477890423784, 0.906698360191899, -5.98655945274833, 2.01695655226225, 
    2.15045238962371, 7.32337061174709, 1.35396093391781, -0.489588429734471, 
    2.72114691086323, 9.44775160448002, -1.09695329052915, 2.65016348203716, 
    3.38145174357922, 5.46239036482249, 7.88387403070818, 0.0462241711403449, 
    -3.36561922488542, 2.58316451070005, 4.7317487616203, -0.285202814929608, 
    3.56559293539597, 5.78587851106226, 4.09472523157281, -0.702924312291116,
  0.119466582555608, -0.366870537856994, 3.15823787419788, 9.396325461396, 
    -2.68266150655204, -1.93237097219506, 0.503818893228463, 
    4.77156199625222, 3.87792511739805, 4.03327416446219, 2.92308693067334, 
    -4.99454020988584, -1.5140579748708, 0.239456657596098, 1.58141412960191, 
    4.93822681405701, 3.47491462919892, -3.45659303589156, 2.83901692928674, 
    3.26844147988861, 3.46432611128899, 5.26141382427486, -2.77861457279793, 
    1.39024722539082, 0.122825353901574, 4.2877322859023, 8.23915181234957, 
    -3.82206196599108, 4.41419253866535, 4.78417682258249, 4.88558485259227, 
    6.59286010972178, -1.45366713877568, -1.81910288722966, 3.56197470706721, 
    6.30248021822672, -2.62812658872139, 4.09391899500015, 9.12718496165533, 
    3.23142378239924,
  -2.15180891507768, 0.390386499261966, 1.73260194170845, 4.57521076326204, 
    3.43273273537056, -3.5451741574528, 0.186954057997641, 
    -0.399576570075182, 4.1405795532443, 8.6072086483714, 4.21543750114098, 
    -0.598674215609964, -2.15656480430327, 3.63172337382171, 
    6.15425194049738, 2.88600407421288, 3.96578679666344, 2.02990558088437, 
    -3.07683578967633, 0.630405714489397, 6.44688271787709, 7.68790117976032, 
    -4.00759035749802, 3.37135780276843, -1.257772499415, 0.476500883774199, 
    4.08948929354927, 6.53834986411965, -4.96696852510896, 0.591880116372553, 
    -1.03129560305596, 0.437316580653459, 3.68744928901864, 6.30874765866533, 
    -3.44946665592879, 0.0966792553747305, 2.62640623295283, 
    9.89419099309568, 1.67944141310633, -0.947240716666506,
  -2.980677406414, 0.930963120535028, 1.05263177742816, 7.22813881631185, 
    4.42888592069847, -4.32640956406172, 1.05152431950126, 6.57117969446264, 
    6.81130112940553, -2.40949567461089, 2.69948377366047, 1.85572846050765, 
    5.65749304602529, 9.04798877841316, 4.52941549892626, 4.73171462538669, 
    3.3279281241325, -2.22850434045128, 0.474708053874749, 0.879160595737821, 
    5.55427800193352, 0.639124244973525, -2.61297641281543, 
    0.603039629489094, 9.52748550558638, 0.618352802146574, 
    -1.14824371262895, -1.87888045460733, 3.30306646649535, 4.1059145234958, 
    -0.836692736248433, 0.861887149859029, 10.5912006569024, 3.3031395555101, 
    -0.243097786710652, 4.66421933456577, 2.45058520423664, 1.73722187186866, 
    3.98137104799937, 4.27901711881189,
  4.5963202770046, 4.54888352477227, 3.41017897530034, 6.98863208816398, 
    3.27272852327572, -4.06126301848802, 2.45247439471624, 7.68707854892746, 
    -1.66974106020946, 2.37057050064795, 3.89013334537838, 8.54098506042944, 
    4.05061687746571, 3.31729989588119, 5.73159197470502, -1.56330916659187, 
    0.404007289173997, 5.67795585253704, 7.56314082187555, 1.42541267995529, 
    3.61985155305146, -0.0485142967857629, -1.27378682842795, 
    1.37265278841456, 6.88511296622361, -3.64071432442621, -2.36009454057943, 
    4.30445534941023, 5.36472856950495, 2.65085743062652, 6.60296316566756, 
    3.64576383470953, 3.51245713937745, 6.00152582611486, 0.626588331720945, 
    -1.44493504086085, 2.37604288854699, 7.51951986302498, 3.76036524192785, 
    -1.20760373010935,
  2.39952516023276, 8.74923047113517, 0.444300992770301, -3.53242579854256, 
    -0.726548692729511, -0.184015263339681, -0.447511793313848, 
    2.60796553450144, 6.19837368947876, -0.619765711949781, 1.99569376592872, 
    10.4080392773198, -0.0909410151147558, 1.45734751786517, 
    5.88107745782803, -0.422657596485724, -1.06939083156885, 
    1.36467773990692, 4.35871705789466, 4.31706865213664, -2.89944683773637, 
    -2.44575702201801, 0.428906424250776, 7.433997931511, 5.36823124250146, 
    -0.588568475992493, -2.30571716153844, 3.37709299382132, 
    4.42032666313833, 4.34426330545153, 8.00069181136796, 1.67740830121304, 
    -6.6979958669983, 0.313530923840976, 6.10118494137149, 9.1870839805614, 
    0.717127742308309, 4.02118321178986, 1.6807986759891, -0.75598777639469,
  0.300209438510171, 5.99934085563491, 1.54742177726074, 0.637405683952943, 
    7.25718985063298, -0.0616302308024066, -3.63671189538536, 
    -1.19996008850765, 8.9130915782717, 2.44729358805807, -3.99411517829009, 
    1.56913302388375, 2.35777418169396, 6.44161132492533, 6.4023963335565, 
    -5.23061710374204, 2.90997395454187, 2.24000883784337, 3.84229856395711, 
    4.23026029516736, 5.06154894003405, 4.17458051341598, -1.3257359909639, 
    -2.11469940670441, 1.54975207740835, 2.36856384679278, 6.55691041710556, 
    -3.75199831260789, -2.88388567500884, -3.31311364977178, 
    4.43699471964038, 3.58602564348173, -2.57248624301608, 2.00117658468557, 
    8.35414146984231, -2.81803833513467, -0.173284127776398, 
    -0.101682478279278, 6.21664535571227, 6.73086036497701,
  5.23463790578384, 9.05023514310895, 1.31925422304151, 0.592913988819645, 
    2.23960232076581, -3.63601889933507, 1.61428661154224, 5.85340391410941, 
    7.8270094449747, 0.442112599896646, -1.95450559958714, 0.668738294110693, 
    1.38969867421304, 3.71870403232779, 5.23797108906815, -4.16664104285475, 
    -0.127633844589448, -2.10246459727372, 6.80425720493802, 
    4.11693534377537, -5.66119105969511, 2.44267493420362, 0.264080319443381, 
    0.460715754067026, 4.11178108759947, 11.4183522346671, 3.91074434046055, 
    2.75413098952192, 6.38861882125533, 0.789437309817596, 0.678085007758019, 
    3.11126364720062, 8.99770533975014, 6.707823043392, -0.0819302179673612, 
    3.8388448433203, 1.45707765164321, -1.51733831233032, 2.2252206873422, 
    3.06545282034143,
  4.84297266828466, 2.89244603255785, -1.83881285000192, 0.201834413638747, 
    5.1281277428912, 4.51352977769236, -1.83187188354763, 1.17946080845811, 
    2.91989187768314, 8.92595453608321, -0.401431574764136, 2.93545897978816, 
    5.22979605793874, 7.76383817547773, 0.0249394928281479, 3.35138337875558, 
    4.54920410905179, 5.14169672178819, 6.26037233334788, 1.53579350949853, 
    0.45330514764564, 5.42587107616317, 6.72524983877267, -5.12432121839709, 
    5.26679091077677, 3.39033144859483, 4.1726848512139, 9.5221286977262, 
    0.504412277533585, 3.56304049966397, 1.14958930361621, 
    -0.442200722824409, 0.290855889651317, 7.3091086922608, 
    -0.0774607801966125, -5.25100041071235, -0.82627819586433, 
    6.32240298759399, 6.79969479190243, -7.31412777025036,
  6.07987724459434, 3.74139468761651, 0.478000961323452, 3.51274403133476, 
    7.7506890936659, -0.964799742453528, 3.69559954219993, 5.41676729521841, 
    8.53479342107432, 2.89709295368997, -1.35663762107201, 7.315405787824, 
    1.91891225083164, -0.704295654355447, 0.177324214081156, 
    7.50205555749565, 6.15000712138855, -1.20097297065024, 3.83220949219484, 
    -0.517672399316451, 1.33215123868865, 2.64179260249043, 6.21678038847529, 
    -2.42188207763828, -5.07228409148774, 0.133156959322138, 
    0.102953667838733, 4.84341394287931, 6.84148699592677, 4.98182931389678, 
    6.05790440727655, 2.27760071402882, -2.67893104955341, 1.43602452735311, 
    6.53816626231686, 2.37717328414989, 0.835601859221129, 4.6896274108875, 
    6.6901475332701, 0.00220939383412824,
  1.24656381872844, 9.03336381194604, 4.48298436049289, 0.670000273540249, 
    2.11788134651129, 0.432112778011075, 4.20553427306006, 7.43544133047633, 
    -2.8907717431681, -0.0326099230519806, 0.913396921308158, 
    2.75143511072714, 7.26448425279, 1.1255696945118, 2.24087417686826, 
    3.51045450186536, 4.38589950846719, 2.64770118305724, -3.40610133450025, 
    1.74557695536853, 2.28288537658426, 7.16158490460563, 3.62425799989544, 
    -6.66284031079122, 1.46464750638271, 6.34092470741758, 0.754523185300485, 
    1.63963738617239, 6.31771831864713, -0.000919603568536972, 
    1.73053143709751, 0.254308038742069, 3.64431868804341, 2.18600899288135, 
    -2.86425027608154, -1.98941087591007, 4.85148009563251, 3.04263903402924, 
    -2.09014328783734, -0.367587865427963,
  2.81829650818446, -2.12827861537559, 0.226955155718439, 3.26946699008878, 
    9.59383817656879, 0.394928079174307, 0.414130497677023, 5.43662717874938, 
    -0.514387080298758, -3.68203819150013, 1.07922137541688, 
    7.28164911375683, 7.82821895548086, 3.05801183461913, -3.09343387643741, 
    1.51142431895311, 5.91277702166423, -1.64894156688308, 1.32221776386271, 
    1.04920658759396, 7.08380976729765, 7.34312154310722, -2.87144914955381, 
    3.43752048254207, 4.5280928008698, -2.47530908425936, 0.698407196713481, 
    -0.0881561099700022, 6.6396740572638, 1.86132891114605, 
    -3.98380295841001, -0.336404676897139, 9.36578753219352, 
    -2.73968126211651, -5.52480143598928, -0.733823573877262, 
    4.95815747885604, 3.32425426666311, 4.14021576652008, 7.5195151488077,
  -2.98763829595963, 1.6114418412019, 4.25093769756929, 7.22492257330048, 
    -1.60557409865748, -3.67844635604049, -0.208888495491835, 
    9.80981372917278, 1.79451846361978, -4.92182278809299, 
    -0.707754548838851, -1.49318547109087, 6.24076921053375, 
    -0.217907608958556, 0.193301347163214, -4.2916111007254, 
    7.10525843448585, 2.41404261701779, -3.33652731686943, 1.41228426494572, 
    1.21847278798029, 6.25771513444638, 2.5294908583823, -1.79572122813639, 
    2.23237201796254, 6.65885662267002, -0.962800510367346, 
    -2.08649622600962, 1.58911331957051, 4.77230366840641, 5.13023250048394, 
    -4.91873637858996, 2.94277173504852, 2.16123521655315, 3.29397266283903, 
    8.11752203752802, 3.48491986124166, 0.381955819892583, 5.01097436148425, 
    1.46329892335051,
  -2.52057088220916, 3.30012224792782, 9.07030064886865, 1.45098019808523, 
    0.773621251750396, -1.43155851492821, -0.842653453439074, 
    9.43692673489456, 3.08584132151334, 1.10938963606312, 6.70444848657871, 
    -1.11983492975046, 0.0539629065232045, -0.633755122002666, 
    3.66938939761706, 9.77684057198918, 2.81258053413902, 5.67722477886921, 
    6.75477886285131, 2.9960015557211, 6.43241816797162, 6.48068703583963, 
    0.983773230701003, 5.93671619979617, 8.91936088975753, -1.12648627440222, 
    0.407570154640851, -1.02990505640109, 0.437603672263037, 9.4653164783232, 
    2.15258744924504, -2.39718827782511, 3.81590988774445, 11.3147625387732, 
    5.63335149407969, 2.59792734809439, 0.89654515090276, -0.291012998329956, 
    5.69555885362767, 2.28889798145782 ;

 tracer_concentration =
  16.5806784755677, 12.8560468218852, 10.0079287795184, 17.7959510273406, 
    14.2147071478427, 18.1146395217204, 18.1055878192977, 16.5752171474429, 
    15.9315284841405, 16.1210578469374, 12.2569383701075, 18.5712427873291, 
    10.2082293224553, 14.2336542378019, 9.42981445143231, 16.360647619035, 
    7.86787390306559, 4.90836851247964, 8.35391862857502, 11.1256412450107, 
    6.8141323736258, 11.4373890843934, 12.0691444845572, 13.9086743886602, 
    12.7401976200924, 10.2934151078779, 8.28828921406116, 8.6662844836562, 
    8.81265948787025, 7.97877252388841, 10.8041720913017, 15.8899314809711, 
    11.2314105053315, 8.26496680938689, 8.87023457704814, 3.60555609856019, 
    14.3353677945604, 7.34489572864561, 11.1068441457843, 9.75843770649823,
  23.7370892359287, 11.6906615102271, 16.2438046383434, 14.1064086235069, 
    16.1494457271729, 11.4314233771159, 14.7360790251113, 15.1283764137043, 
    12.9805859824249, 7.20752933949203, 11.3572514733244, 2.85732820323162, 
    8.93997198301381, 10.1991999982648, 6.36206547526902, 8.25641307132968, 
    3.21793770162348, 1.16170652079105, 2.15615282527821, -0.449761102212168, 
    0.466738649171873, 8.4314889403394, 7.69877045253646, 11.2273580402091, 
    9.32869425323132, 12.0068383536231, 17.9648000722638, 16.3638950560236, 
    15.4536129544142, 18.930551244709, 18.7893930554259, 14.5475600185335, 
    12.3464007951362, 13.5324283550188, 11.263437020787, 10.750984036141, 
    16.6468336220236, 18.1711928176268, 17.5823322535446, 16.2479368017635,
  18.7910713857628, 10.1885474659741, 10.683327618907, 15.2639743019514, 
    9.54975607443627, 10.6095062592655, 8.73275604601887, 11.3197801971763, 
    8.84938259465884, 8.28617201516776, 8.50909567576895, 5.85228778528183, 
    12.2351576891107, 9.52499150677607, 12.1552827465839, 14.707014896531, 
    11.5366125242202, 6.12148142099447, 10.7634162370086, 7.49196015860538, 
    6.51386869731791, 9.04394132587517, 11.9619040491267, 15.6269250433156, 
    8.95108711480148, 9.76091900528363, 13.5677716841454, 14.6672836769504, 
    12.8467621984957, 8.83283902146145, 14.0996978507217, 9.98460066096133, 
    7.4631225791385, 11.0826659094975, 8.76405397530142, 8.02414782609398, 
    17.3264939872335, 14.503168647341, 16.6445854731839, 10.0635669404357,
  2.77498230888648, 8.44571730064523, -4.1197343130417, -3.06214786003408, 
    3.22779378212245, -5.47782597857801, -0.426271363444418, 
    -2.21437765855779, 0.0111112098948758, 1.17608807121593, 
    -0.337770223615034, 0.461816953648062, -5.58931671766332, 
    -1.78671470906829, -1.04326492107822, -3.22237278600678, 
    -4.08536266660411, -6.03078054640007, -7.4137775204439, 
    -4.45012787861488, -3.06181689221031, -5.89216540639877, 
    -6.29958114133866, -5.83665372824471, -5.96131249708971, 
    -5.33750197000785, -0.165583372587333, 1.40158688179315, 
    0.121029078450554, 0.454225283111805, 3.15598590762142, 4.07622044774769, 
    1.41259373085383, 2.11029513336322, 1.67420666563757, 3.75792011113633, 
    -0.160857761121339, -2.84592216157862, -4.3846808248899, 
    -0.618160028970105,
  19.4681691837424, 25.2897100216978, 25.4785932465922, 26.4921805403799, 
    25.0429870282825, 26.5546107497891, 21.2609641687739, 19.9002127557462, 
    17.247973303896, 18.9420569689686, 16.0446185704737, 15.9737954256288, 
    13.4731494491713, 17.7971904492463, 16.4682892893815, 11.4997298787808, 
    10.4052788193488, 8.03773146725062, 15.0206464628892, 6.89915327546297, 
    8.70535573447495, 4.50947974228785, 9.74763384334258, 2.275969575996, 
    -5.82656148988758, -2.72791451790695, 0.638933616334362, 
    -3.40352428224385, 1.43607008099097, 2.64153476459198, 6.11259281868653, 
    -2.86748944518192, 0.823217470140268, 3.81121166211183, 5.37611559127017, 
    4.61321553268875, 12.6131805502779, 10.6528672514774, 12.6982645801609, 
    9.63243245170008,
  21.58906768641, 16.5799537652425, 12.3086825725434, 13.752106421104, 
    9.64034926158402, 13.8311131029561, 15.575080938664, 12.442831352054, 
    14.5613038082586, 18.3546084019746, 18.3694342334502, 18.5014417144717, 
    25.1817884347161, 19.5194358017226, 23.5648824158626, 22.2789065475322, 
    21.8473861537678, 22.4550631241139, 21.2638612168639, 25.6897356001354, 
    25.1336318470598, 32.7164253595191, 26.8134456972647, 26.4249133077711, 
    23.0366460321926, 23.718183715109, 21.484081010722, 20.4436042204872, 
    16.3388845231938, 18.052612360683, 13.0547289907817, 20.9218273440486, 
    17.6734956871944, 19.583903798883, 22.4514012112422, 18.5904363908674, 
    12.5393039589467, 12.7731935675803, 13.2324587308347, 7.15690753137431,
  -6.02968124290731, -0.964129903517134, -2.52269513604177, 
    -1.05453358049688, -2.22605136573904, -3.75757327740113, 
    1.62149487343458, -1.16975386653792, -1.084779521611, -0.139989592695651, 
    -2.77247152972151, -3.54755282863257, -9.30571041872541, 
    -5.47180728831169, -8.2967109371731, -6.29848547854908, 
    -8.45805700718076, -11.6045979590215, -14.1925999098826, 
    -12.2962747511491, -15.981699130033, -12.396038993146, -16.5533733281545, 
    -14.4252053430503, -10.2862549926317, -16.2337997803208, 
    -10.5880618585974, -13.3886066453468, -16.7222406210643, 
    -14.3420087329354, -15.46364265479, -15.4679619600513, -15.8152210466875, 
    -13.221466238895, -13.9569013992442, -14.3444777153192, 
    -12.7368490024893, 10.2104568738866, -9.19622341899567, 5.26406606095984,
  11.2671810594023, 7.28966170168189, 2.59968964618431, 7.75703759216458, 
    4.73109897877386, 7.99764302054806, 7.12114019163135, 4.25417859917641, 
    4.2708735550596, 6.93268657889847, 1.36444753907404, 3.80867021493252, 
    3.87251232400103, 5.99895059647915, 6.16865788534952, 6.82753810683251, 
    0.593164258219324, -1.23202528631448, -0.458160891016947, 
    2.28049042841114, 2.54225406447941, 2.36706150654672, 5.09873933180906, 
    4.51292880187263, 2.86266783572437, 7.33397375287864, 2.77790643482202, 
    -1.79328301159176, -7.57815716553773, -2.67947730902001, 
    -8.65145403520214, -4.49230566128944, -6.54302716417171, 
    -1.98541725719021, 16.8339359098169, 2.91298007720121, 15.7881917693899, 
    3.05271803079137, 8.17006157632624, 4.05219124847325,
  24.9780802704011, 25.0403011836274, 23.392234531611, 25.1628151674873, 
    20.3565276610036, 20.1325538935175, 17.5057667879394, 19.9717861052116, 
    15.1336233803121, 13.8157242504443, 11.5848275721075, 16.8985080073793, 
    16.2668286756624, 13.0944142858267, 15.0769426795788, 5.1019579781365, 
    10.5513254343654, 9.95023310904584, 15.5085302530333, 17.7878006134904, 
    14.6124694406347, 17.4235706988286, 22.7190936235718, 21.6320605918898, 
    20.8107873532909, 23.0245391969157, 24.7108308178843, 22.1198334850662, 
    24.5445808096252, 24.570234812068, 26.7515050215498, 20.6167319001511, 
    22.0590031039811, 23.9068484256057, 20.8743362833782, 21.7871375809374, 
    19.7953260335811, 22.2769673523468, 16.928774030199, 16.5854093319081,
  -1.71100484721205, -4.18804131838736, -4.79020245357755, -2.80870862837262, 
    -2.41530842022608, 3.09843169919832, -0.51201186971613, 1.95094933634979, 
    0.122503385950321, 2.7563984058041, -0.911559855339908, 
    -2.54750231259306, 0.305073903341739, 0.108173765779973, 
    -3.72277390891085, -3.298807675439, -2.94241034136695, -1.04631654894691, 
    -4.40272340304488, -4.89643869899906, -1.0328432592063, 
    -4.49989752988113, -4.26627356943548, -5.29365248921276, 
    0.102953516454976, 3.4587678722946, 2.65872821870641, -7.7961517732276, 
    -2.55649987354911, -2.41760362891413, -4.68519136213278, 
    -4.05813737348734, -5.9462546045169, -7.09722117722918, 
    -6.18870704481811, -3.8459660113255, -2.0537684764472, 1.34346895219315, 
    -4.37952637124473, -0.493974096436032,
  -4.42050893719967, -5.50034278864229, -2.96512954027901, -7.44319905139082, 
    -10.4614668442621, -8.87549994683128, -9.85269804749553, 
    -11.9293544657532, -12.5650945101882, -13.3163411018152, 
    -11.0706049292762, -13.0114923730998, -4.99422551362893, 
    -13.7164523734475, -2.01866202036612, 0.782044304446279, 
    1.09185858829763, -1.947454271048, 0.731296680757365, 1.08129295046847, 
    0.378095256982842, -1.33642624781946, 0.341678473334423, 
    -2.09801421399728, -1.85146360977758, -4.44822213746556, 
    0.791766741113215, -1.44420615264729, -5.20529505429213, 
    -2.63744842792202, -7.87654812449424, -4.47665762582176, 
    -8.68475433961269, -4.24723532332229, -9.80169699354551, 
    1.61454466253905, -3.16435757529997, -6.72049230419065, -8.3557448373307, 
    -10.4179505455966,
  8.77742018258262, 3.46348083490902, 2.56438792792127, 3.43402397818483, 
    5.71638452697153, 9.50878105541744, 6.12771916687423, 16.9994082233618, 
    13.4558613216982, 13.2836757480142, 16.1133438024988, 14.163490629551, 
    12.9024085072314, 12.5958647681168, 14.5827297431564, 9.86089466132964, 
    13.57913755745, -4.02150231858522, 12.7824467418575, 17.7233747010498, 
    -5.06110672664498, 5.24865885958875, 1.49765299552606, 2.3628690099947, 
    -1.19445439476253, 5.42445881158401, -1.58422118997504, 1.15428555752381, 
    8.25130031595351, 8.61754821612098, 6.17316092590757, 9.37516773378483, 
    7.92754839727775, 9.16937347516802, 4.3260118550599, 3.7997428045899, 
    5.15041545135845, 4.36881707456634, 4.00979113387558, 2.63666310323569,
  6.47783801529701, 2.30044821888948, 4.13710638678479, 5.15464287670356, 
    4.02564407187907, 4.53059380973797, 5.45079148494393, 2.25303063098438, 
    5.77468464890538, 9.92620640634305, 11.6233946914202, 6.98271383095647, 
    8.7539728559947, 5.66978953909201, 3.46441752491621, 3.367732113292, 
    3.17968939808208, 0.89993407888152, 6.84860734893927, 8.86569760399324, 
    7.88453976412414, 5.23993863008684, 8.44775417656553, 2.8254896099347, 
    7.0745651012811, 11.0282938882699, 12.1072866723759, 16.8522335272203, 
    8.78402162958169, 16.1816876228875, 9.10783778928691, 8.38411626030058, 
    14.6039976884715, 7.6967603613587, 5.2687014829145, 7.1799562482178, 
    5.10320835592947, 3.51360206455203, 0.657981317434688, 4.10551298813819,
  8.42139319818166, 10.0812637760885, 4.84606826683333, 0.262796055722062, 
    2.19838140173279, 1.42530636482948, -3.57390585369655, -1.80618894286937, 
    -4.52590257274401, 0.627097813041243, 3.34466093814858, 
    -6.02894508567305, -4.57505114529052, -2.61710558238829, 
    -6.45540678482208, -6.07362872613641, -2.11839608115887, 
    -8.59404341711687, -6.1629256167998, -2.12385520167636, 
    -1.93047788525158, 0.0106843189382142, -0.54251954713786, 
    12.2492815162848, 13.8904263502053, 9.02719509768859, 8.84543996348015, 
    4.69557847269975, 5.83207233558566, 7.83736127578551, 12.3412925388182, 
    10.6990044048318, 9.76995315848689, 7.22407522408253, 6.59930977756965, 
    2.18432366572923, 4.88873157343505, 2.97462861859745, 7.45452561763432, 
    3.94243188508147,
  3.53535098978011, 3.11255618765266, 3.66443712012932, 6.10600602635868, 
    9.63596866037289, 9.19342391494896, 10.1867965764653, 8.57168290032839, 
    10.1995939419086, 13.1152553446255, 7.33909434350162, 9.95620841602496, 
    10.1692463023613, 12.6026045718287, 16.5800010537689, 13.2022304890196, 
    17.5952324460914, 15.8681454995441, 15.7377284268499, 14.7401543601497, 
    15.0671689099872, 13.573591974561, 13.5677463771767, 13.3173569322172, 
    9.2088276560324, 11.6500881781987, 11.2283634216955, 10.7213847494202, 
    6.72147381752761, 6.6740880668788, 6.5010081798936, 5.88388747141236, 
    6.18950769118055, 6.75693966357353, 11.3577496978932, 3.78618090994803, 
    -3.4373388497125, 9.48920234430454, -1.8422892122503, 4.59786393516717,
  13.7762260714692, 7.50214541217701, 12.0309439894463, 9.00820040654582, 
    4.9621109023979, 4.15667552696578, 3.57551594716883, 2.62590886887841, 
    0.738444822887616, 4.75944878445406, 0.365150754724155, 17.5759406998132, 
    15.0142109945543, 17.2330740879274, 8.00095038968608, 11.1467952250433, 
    10.5409347559468, 17.5124649643856, 12.5427519989923, 12.1571420571219, 
    12.3876271486183, 8.16565144489264, 9.11144237594664, 11.2027226359733, 
    8.83786516361147, 4.80497219708305, 7.67398769042229, 7.32098620239909, 
    3.23539007042195, 7.13276561857565, 8.38546415559468, 10.3992392952375, 
    6.32758658582085, 9.9123090820992, 7.50045442950832, 8.85488473608179, 
    11.4670785423877, 8.1181976065651, 7.14239427846599, 6.22306845752127,
  -4.98925073869639, -10.143161162952, -7.44042682276071, -8.79400795083691, 
    -3.16984312468101, -10.8465077789636, -8.37222531901539, 
    -12.5728515352332, -8.53904245470682, -7.74782188419016, 
    -8.86353243440369, -10.5070952426966, -9.88591326166695, 
    -8.04818446063482, -8.94735729287236, -6.97128270340959, 
    -7.68023823680485, -7.9515530907139, -11.431889751859, -11.3332694448768, 
    -11.6825274462174, -8.83021529727189, -8.92942915730616, 
    -9.37959166482097, -4.63878373408957, -4.63439965897814, 
    -10.273302767786, -8.31356372933308, -6.2525277346977, -11.1800829322018, 
    -11.3577727588517, -13.9982316086236, -14.5583750854268, 
    -13.1985605943372, -13.553308707562, -15.1739927775769, 
    -9.14876364918448, -14.5274756489619, -11.6331921171252, -8.85549333964233,
  12.1240781210244, 7.53568803398636, 1.55803536417351, 8.42959793641696, 
    3.01531957486193, 3.3731000585926, 8.34179768502084, 7.94260980480812, 
    11.5546116853466, 6.89275286837712, 14.8106988350073, 10.9902159377046, 
    12.9049163300148, 12.8868666455111, 10.3077131952403, 9.84220521828877, 
    11.8657804927762, 7.76374877785249, 10.0614593430303, 12.8081590367362, 
    11.0401178059154, 17.8123493140266, 18.0947767535728, 14.7035306727019, 
    12.2928615960656, 11.0982426664841, 11.7719606448948, 15.2624971727029, 
    12.9207839058306, 14.6690200057039, 10.6926427557888, 12.0645185250548, 
    10.5012688759799, 6.07210637080156, 7.28792334905541, 2.98000452596735, 
    9.20798373326447, 6.32883447974558, 9.02054075998598, 6.91971211348219,
  12.1777414664911, -3.03911517502881, -4.15826596040283, 13.0733164619758, 
    -4.70022833231206, 1.15649886728931, -4.51253697355867, 1.5007857166132, 
    -0.9299501666105, 0.891676475886141, 12.0153548911527, 6.77926678773399, 
    2.86730185066516, -2.31003007243998, -2.1048602426959, -7.04276108787679, 
    -12.6027514779369, -9.20902322050914, -3.24729923005294, 
    -8.34064416790766, -3.53247984375765, -1.90831583966701, 
    -5.67032807056763, -1.71100034423886, -2.31065113229713, 
    -6.51318982304097, 7.8674215225239, -10.2584780844692, 
    -0.208923814333723, -11.2308378401002, -9.83259798878648, 
    -6.67764078221564, -15.329947345633, -3.1141624368166, -8.62008674328647, 
    -6.29056243740714, -8.48478299096418, -8.92313144275965, 
    -14.4021418156017, -5.90623383816503,
  12.3852984262078, 6.48365660567171, 13.498680703859, 8.92108256062539, 
    14.0077503396671, 14.5000156423473, 12.1209292477521, 14.4779365012879, 
    20.4968360839585, 15.0898576092638, 22.4754998514491, 22.5361153352184, 
    17.9311554716297, 31.5869626852565, 23.2793061182168, 25.8129676596798, 
    29.6732409554888, 29.4741226333835, 28.618194394406, 20.8547318218684, 
    29.2840553660311, 23.2206098500631, 21.1881405523818, 21.0942016311974, 
    17.8792128863295, 22.8197441564074, 31.2307597084292, 29.9797805365049, 
    23.9554075988684, 28.0907699782973, 27.6141563135366, 21.1022428936917, 
    19.2270403776051, 13.7951617495471, 14.5359764226152, 14.3926439381165, 
    10.8101099663907, 13.9757290095602, 8.28216800455389, 10.4952481104216,
  17.8181102691507, 24.5405182841117, 22.2366502613092, 18.916386475505, 
    18.7314764185495, 23.5232596331651, 26.8615943846296, 0.535941979495145, 
    17.3245687852843, -1.7531359768382, 7.73424231863811, 13.9049326954119, 
    9.40136920796423, 11.6657246744534, 8.23369447786012, 6.2535900781065, 
    5.72982853891686, 12.7750544633643, 6.15709072397456, 0.414239164015562, 
    3.14663040638352, -0.125766042164567, 3.77907957707374, 5.7177140747615, 
    1.96636533766954, 5.95593627397898, 5.95402472354063, 4.99048139746362, 
    4.81155907549732, 5.67879564441908, 5.60062363641944, 13.6202185720188, 
    14.741787332634, 12.515836004341, 9.14539575387398, 14.1745933546396, 
    12.9599704594654, 12.5073080070653, 11.7539481594278, 13.9747294373645,
  7.38442803134356, 4.57293624614997, 7.87344637881972, 4.7843952972277, 
    2.45074490137687, 6.92423539075071, 3.19957095761173, 8.96111097708558, 
    3.9135892586066, 1.01710081351429, 7.4665073511655, 7.45377525168753, 
    1.70939661585804, 5.15214955072529, 9.43932077651803, 13.0557067808155, 
    10.2264483224886, 12.7963393424842, 13.2937320215668, 10.8266738862537, 
    12.0980786569754, 8.39918096676942, 10.7708175920641, 8.42838112074727, 
    9.04546371605483, 7.75442714641856, 6.52365558943782, 4.46197718529445, 
    4.08618582475488, 4.02917138741194, -0.501541213547934, 1.31258532300574, 
    4.35713286367203, -1.78985224113237, 0.843308848905569, 1.73223766431291, 
    0.0534451697074058, 1.94639267930318, 2.01025783086159, 2.77283112238832,
  -6.75213157533525, -4.22146547217889, -1.89510472494074, -5.05321469587411, 
    -5.52858133595581, -7.42000416899467, -5.24199509837469, 
    -7.09406811024661, -8.37950018943844, -6.71640807521146, 
    -17.2995696791913, -19.1818300092793, -9.9113490916178, 
    -17.9079305851684, -28.1386350742491, -14.5000771333996, 
    -17.3579000219336, -17.0918170359846, -13.4317701690791, 
    -20.0196018324913, -18.2720409531746, -12.3937120801341, 
    -16.2821219781051, -16.5602794364633, -14.544395451021, 
    -15.3495374085187, -7.06993513938499, -12.7610965560076, 
    -9.90976868966766, -7.38687024233682, -9.91315283073756, 
    -7.30122619223603, -0.724470551714198, 0.764596020478353, 
    -2.83462028623025, -1.90275085462086, -1.07884523777618, 
    3.33047502064932, -19.1698939495127, 2.5946604846875,
  23.1118226284658, 20.8282206836571, 23.2871069914039, 22.1567843848576, 
    23.4846265752984, 22.5566783082877, 27.2568887096182, 24.1872425694866, 
    13.4644873820782, 19.3983622637527, 16.4086680688316, 20.6119570225076, 
    18.8180568225543, 23.2747139761553, 22.0638844185218, 21.2020433085993, 
    16.205009070075, 0.943078372589839, 16.5616671817646, 6.94106363866284, 
    10.8092172732155, 3.40998775498038, 2.86782371096762, 6.22987212948406, 
    11.4181446367194, 8.75051070242346, 15.320017848632, 14.505885717998, 
    16.107894860373, 17.6733090255957, 20.4263011677002, 17.0020771928123, 
    25.003291790433, 15.2070349420429, 17.0867328671628, 21.6682944699099, 
    15.3713578450101, 22.0992297576825, 17.6236463680907, 20.0217756641596,
  -4.52138086332201, -13.4343494136374, -8.33318451214252, -9.11286492175584, 
    -7.55230444247097, -10.719148532996, -10.162791396556, 3.0167931462575, 
    -10.1443126483926, -6.939135108563, -3.76418680457489, -6.78617568469299, 
    -3.8191680756336, -4.63720292440145, -7.79435454830203, 
    -11.3689885359119, -7.17816199921805, -12.9584658130826, 
    -15.6575763240267, -11.840395458069, -12.8389274700686, 
    -11.2002995740487, -12.3418632114821, -11.773492653408, 
    -6.67128995105491, -6.73210376192438, -8.452503363406, -10.3396868876665, 
    -14.9096800172948, 4.32338758834979, 4.79660928583878, 5.86170100749943, 
    5.96456547624949, 2.97253898788931, 2.80279824993083, 3.57110901094728, 
    1.9777691878512, 2.7353709100994, -14.0501372487744, -3.65055603649476,
  8.46117565329877, 3.29597207955531, 3.66279573304536, -6.62315295250721, 
    4.90304578201303, 2.49686191353234, 6.65953022608952, 3.82663762434737, 
    1.39985025401191, -2.92667702846639, -0.775192052958899, 
    1.61185229480264, 1.90225089407365, -0.699701196589021, 
    -0.572305845520399, 2.25548643086705, -1.96430073181917, 
    -2.70857552340189, -0.763629045052462, -5.47306774042419, 
    -0.355325776796977, 1.78156650510355, -4.05765825388494, 
    -0.772910080241913, 0.918559973820588, -2.81576254035061, 
    -3.2361999714582, -0.974917164280434, -2.78318191015937, 
    -1.25372775569797, -1.77532217691091, 2.30056811157366, 
    -1.44233965832957, 3.54749032164993, 1.45555115033705, 5.04135943952458, 
    3.09046010348682, 7.01972619392702, 2.24870093855281, 6.93357837218224,
  22.4746935458122, -3.29269074388963, 19.1060171687199, 7.86110516055374, 
    4.78022937035865, 18.750413002954, 6.81187389921344, 5.81097904081213, 
    6.5119595893928, 3.5867017168073, -2.83278709720418, -2.5333315174624, 
    0.750731507391088, -3.34960665139649, -1.91271206033684, 
    -1.93335200537824, -3.38400983479647, -1.2726297785999, 2.99198537402597, 
    -0.283474974859548, -2.76129267627936, 1.16900760222607, 
    -5.20277469325713, -3.77120364271111, -6.39152331039015, 
    -3.11486207075432, -3.06342343781646, -2.7162155516841, 
    0.144672264474073, 2.47739243657558, 3.56060754480274, 4.57705094185092, 
    6.20278437732522, 3.74261894827907, 3.45246641743393, 0.971482623555017, 
    -0.353783299987546, -1.9095417605932, 0.144718393689897, 1.77679413463276,
  12.0755191939227, 14.793909313518, 12.7859885491631, 8.38504930182929, 
    12.9193894479023, 7.1733739776557, 7.42413187164554, 9.58745539570773, 
    7.60903197001914, 10.9241426765319, 11.2065630942921, 10.4443377230791, 
    12.4272783739695, 8.99693289243366, 13.6837768030301, 5.19464497817844, 
    8.75212525089863, 5.04622812503167, 9.98095490586331, 4.01369524777643, 
    8.67012991015134, 7.58962727909053, 10.220584340582, 11.6468243252448, 
    10.5530622618738, 15.0172306502654, 11.8393153148398, 13.8079354709662, 
    14.8333036863571, 11.3584723213133, 15.2477878409664, 15.1168800680108, 
    16.1296962787346, 7.98495401093875, 16.6441127854455, 11.7336251782221, 
    9.04250185770656, 11.4907472662386, 7.15524943489465, 7.80453325163253,
  -2.35022579363419, -6.829235590064, -2.216486614012, 0.596997052689681, 
    -5.53021578493478, -7.66591812474922, -5.01131410969628, 
    -2.60846332114872, 0.334356999551745, -4.88517214982644, 
    -0.0413926550383348, 2.49096222078172, 5.74177982155809, 3.4825268968392, 
    2.15305994436244, -1.29335044178201, 5.00556514079838, 0.332848547927349, 
    -4.49743239624353, -4.03977580407696, -2.86738655937675, 
    -4.6184609579464, -4.51355069681209, -9.03366913008622, 
    -9.34588092285128, -8.64235155900702, -8.68827019637655, 
    -6.72835007537209, -4.96317556312484, -8.26204238775829, 
    -15.4218879185069, -15.329193967467, -17.8337510869503, 
    -15.1481863272281, -16.4778575322296, -17.8057819702525, 
    -15.6611175092283, -13.2933841090627, -18.9590808182099, -16.7340401230137,
  18.206770657028, 13.5777193208487, 17.616794629567, 15.4955737004995, 
    17.0584415937586, 8.88782745908963, 12.5204913989301, 12.6070944501761, 
    8.82905022191161, 7.4205648262138, 8.14499994435887, 4.74513463921521, 
    7.66231188128256, 6.55815222529207, 6.0520895690216, 7.75180069836903, 
    3.59470971215228, 5.97731673464396, 1.94984518877916, 5.09054890667142, 
    4.48456752877349, 6.03626120600721, 2.75534757851812, 3.37506752112456, 
    6.73663064283013, 7.226840405823, 6.02286833690356, 2.74280986832281, 
    5.87094318248816, -0.715363474968128, 1.9084330886375, -2.99995765059446, 
    4.06749968040746, 4.00158174944131, 5.85111003772316, 6.43969708246546, 
    0.776144531460645, 1.19918565990815, 0.493258234272806, 5.12076906418084,
  -0.253254105637225, -0.879131431323352, -2.19063091230455, 
    3.57594754098591, -1.11568043653472, 1.88049465009402, 2.04138864554183, 
    1.99011805693335, 2.07228490081825, 0.561978978206044, 
    -0.738019655808289, 2.83612533962207, 5.60032740012733, 2.45734945304583, 
    7.73612790269865, 10.081351937788, 13.3335163400982, 10.8277728387109, 
    10.6653650286831, 12.4715399998752, 9.37962346404347, 12.565979296973, 
    9.30511462341618, 14.0660818902846, 9.85320555768432, 6.44002695156067, 
    -7.90823477852657, 3.91296798801453, -6.09765281988378, 
    0.771301195539059, 0.466575364670471, 0.19915945333298, 
    -5.50048665475737, 4.02952980795651, -4.09863025031997, 
    -5.81369421868192, -5.28520143960182, -6.60286859325054, 
    -5.91946222557075, -3.02144637592728,
  11.9372242595181, 3.81123521223507, 14.1117722355567, 10.8516312502803, 
    11.2384489564935, 11.7386845951427, 14.99844493192, 16.1389802834219, 
    14.638547889108, 14.7347671504701, 12.6486792930058, 16.7086673863952, 
    11.9882504162757, 15.1010570116034, 15.0473663658799, 13.093135053748, 
    14.1596200795189, 11.9735012366605, 14.3852266058255, 11.2751435392616, 
    7.60386356328515, -1.78164586125143, -0.986660072081292, 
    10.7315463665636, 2.59551865579955, 6.45040317360358, -0.382301669958925, 
    4.38883906404189, 0.237995308175766, 4.97402156772567, 2.16566110114101, 
    4.96461569437602, -1.03078321222777, -0.306366213442638, 
    4.91884515202968, 3.53964326067077, -0.739881247672235, 
    -3.70038222311589, -0.773894481545014, 0.0933985441149659,
  10.1841320544014, 4.72333574652061, 6.33909477007974, 3.2528686935872, 
    3.93989617611355, 3.81858591875306, -5.54836398080405, -1.20833219189757, 
    3.18850871851124, 1.07782417037489, 6.222265423225, 2.54375535369207, 
    2.12391992998975, 5.29157108352372, 3.82568848459465, 5.14873500962078, 
    1.00312565826949, 3.34079690238931, 3.74248669966198, 4.0305694887943, 
    2.1592809107256, 0.671533322318702, 1.68062817597573, 6.02999943092375, 
    4.69808148736737, 5.90133070055372, 9.08829718401073, 9.53365763048556, 
    16.2452419972544, 13.7829856257118, 11.6239521150072, 12.1052276139151, 
    2.79881069774935, 3.24715315956509, 10.6027933824411, 5.28009308016806, 
    8.33815007511991, 3.16709013694113, 8.55163812002153, 9.30283793110462,
  5.57122072050014, 5.12896958614946, 2.09051390775165, -1.32614078633215, 
    3.10371259091032, 10.2658920648013, 8.46709704344097, 10.384300603859, 
    11.40186604613, 9.53574511224688, 13.6441378498548, 11.3787136335365, 
    13.9535333890184, 12.8214620372344, 13.3768776524961, 8.78087053995151, 
    17.2063244659519, 24.6339899704751, 6.8755340583884, 24.5512285971183, 
    21.7319926567959, 24.6157885358805, 20.745408920434, 12.6324318075817, 
    11.0570786575786, 17.503136458669, 7.58816909232527, 3.82110432118067, 
    8.10303940856043, 7.83501043347261, 7.76606965172855, 8.86485772340061, 
    8.26046046334805, 6.2782701745633, 2.83611914590421, 10.0583769796592, 
    5.65094820697277, 4.98024483063696, 6.7125783758448, 5.19032184922014,
  0.393291616441586, 4.94326065878336, 7.63650486038094, 8.57162353252139, 
    7.36028543295989, 10.5942914030695, 13.497103580181, 10.4895013968373, 
    8.35114848686257, 12.0676498384293, 8.22001914580983, 12.3277656787754, 
    4.63740490571034, 3.88954494259333, 4.33510520474184, 1.94862596614512, 
    3.09511963431775, 1.72268655575307, 1.99208225442809, 4.78046703904022, 
    2.00114796406448, 4.64168122837501, 5.8616798313344, -4.96184156526128, 
    5.00927333561458, 0.912114221017771, 1.39889617097742, -5.27082082281545, 
    0.0186457923027467, -6.21089184867173, 1.64651927230812, 
    -0.861569556875528, 0.09281146475849, 5.18710635852085, 2.13169181095507, 
    3.5188835131243, 2.51020709398113, 1.10385714118743, -0.106396380629136, 
    3.79828507706885,
  14.6480099920471, 4.55012646439504, 7.6627896958481, 0.847730497509377, 
    5.2292040880598, 6.07838069942434, 4.90343495180711, 3.19840632332681, 
    1.80234298180698, 1.37996088916566, 3.11539643724254, 0.13431046373562, 
    4.61414273590975, 4.30941600585028, 5.24517763394115, 8.24973859988, 
    -1.30321423150085, -0.372089555777458, -4.93633559018195, 
    -4.56866560767005, -0.610812089265747, -5.29318223479298, 
    -1.54664309501362, 2.02915188215177, 19.2765766019175, 18.7820786044945, 
    16.1081424169931, 20.9760360743237, 18.0205206328341, 15.1542706024574, 
    21.5944353091039, 15.8519829394771, 7.05120340499577, 15.1753578303753, 
    10.3835690186216, 11.2439716521586, 6.7447827904316, 8.66517402133851, 
    12.5014092395692, 11.5962124523549,
  18.8622850592421, 12.5651391190344, 15.889851126772, 15.4869042186963, 
    17.6971591473443, 19.0833347499578, 18.1666275208721, 14.8736205200765, 
    11.8538267789872, 14.2920755401803, 15.5377646769452, 14.0398370609732, 
    12.9368853755723, 10.1959837717459, 14.5842358617433, 10.5556101352032, 
    11.9154766996096, 9.68334559299747, 8.71648702609506, 8.81402656937017, 
    9.3018489742844, 5.25702229455882, 9.55215620733277, 9.20271253503598, 
    7.21500147231723, 8.03012749963699, 5.21449770474042, 8.65970849690898, 
    7.81356281203781, 7.62864721138039, 6.66496175413379, 6.58500585412567, 
    5.21278922218792, 11.4914170853353, 15.9078835353261, 11.0089250205124, 
    15.1096555324108, 12.9280334309382, 14.6105107420691, 12.0780812090979,
  0.910845854424799, 5.09169167406427, 4.33839883139241, 4.51320096466423, 
    2.10845036651298, -2.84045072910295, -3.42220272451146, 
    -1.87627505779157, -5.21112539204646, -27.4888266847458, 
    -10.2522181241014, -4.36634859372666, -27.5548347931698, 
    -8.50136639937224, -20.5165371589311, -16.3205873951774, 
    -11.1900920123601, -18.0466656334256, -14.2942078598055, 
    -13.0142167076848, -18.8857333786585, -16.9931625874155, 
    -8.83720983505131, -19.1158384916744, -10.2973279432687, 
    -5.70679245401279, -6.2120911653635, -5.76200889511063, 
    -4.03900425503765, -6.64439797326184, 1.97090275313213, 
    -3.02071421969392, -1.94640738300108, -4.90892346353444, 
    -8.49388935333239, -10.6517523878133, -7.58711895513539, 
    -6.34579462110507, -5.4541659843749, -7.26999994067962,
  9.73132397662618, -1.44421112797067, 6.70445659036644, 6.74739065174997, 
    5.75831184347716, -3.01145086243488, -2.63418377830128, 4.3760024504086, 
    -3.71855933409463, -5.26363832534697, -6.86444836672284, 
    -7.02732290440961, -7.02427663746455, -6.08464781680355, 
    -7.62734248732387, -5.51930400978842, -1.01935439710213, 
    -3.26509627302652, -5.4429437758809, -2.11950986874791, 
    -5.88027408725402, -1.84883526596029, -5.84760471605238, 
    -1.9910812512926, -8.1664373150004, -5.05597630650749, -6.62844542012747, 
    -4.08920410711694, -5.03841617355682, -7.12687032373524, 
    -4.05063257549139, -6.03970041865169, -2.66425883599502, -3.829011648127, 
    -3.73069987558696, -4.44845975714719, -2.38191659146699, 
    -1.96911721420413, 1.5099587647845, 0.772567116712742,
  0.674897204605106, -5.37551062735477, -11.2586155028753, -6.56955273989126, 
    -11.3227129428136, -5.13473339201743, -1.78097664633226, 
    -4.86644634852279, 0.923675901693596, -0.240852390249431, 
    -1.5316549679894, -3.09807824458031, -2.65998089764366, 
    -3.74783278187556, -0.910330031981113, -1.3405514430352, 
    2.45006286415247, 0.744317342781487, 4.2614681497258, 1.20527264213814, 
    3.00013090148616, 6.99897066603118, 6.21300394998094, 4.41809628949404, 
    8.18068162828988, 3.77715752235431, -1.50394439065358, 0.882395659432233, 
    2.40187761547805, -2.21719464553263, 0.251353037077164, 1.04658937746775, 
    -0.464584323071585, -4.47111584372381, 2.03585810658903, 
    -3.12195249413281, -0.600435242437765, -1.9762367199066, 
    -5.03091011389575, -5.89928089851793 ;

 source =
  107.570750308843, 15.8229757542169, 15.5467186048927, 88.4739611364023, 
    22.5671250146668, 74.790002832312, 86.9660699437604, 44.3902416261048, 
    -18.4703719137213, -9.30913972931679, -75.2491813660742, 
    80.9353984035727, -106.382091363384, 38.2686838421412, -5.01032047802736, 
    76.7078146607153, -105.763708784661, -42.6727773932221, 25.2573567270154, 
    1.70668200899826, -3.61802911862134, -4.8707681180841, 25.9203928692918, 
    60.7403605066034, 63.9208932211252, -50.6830393787446, -40.4541633641759, 
    -10.8323386994894, -1.69693924446176, -20.0412871594697, 
    40.2987170080281, 73.1754441355168, -5.49292437738618, 1.09479652699369, 
    9.10620784368974, -101.903986027355, 115.924876510301, 6.22873299125757, 
    31.0522935221909, -42.2119766766289,
  177.138228061098, -20.3771229164499, -41.4199386618604, 51.9703900414156, 
    4.08750677323563, -36.0094902742802, -30.9840531480087, 
    -20.1997197351106, -31.1639412621739, -7.49558898724971, 
    41.1913647577225, -66.1253148744295, 1.86439483405112, 48.5405382402888, 
    -2.84639423442412, 7.4970836522742, -59.0460314101673, -45.5596993851044, 
    2.78817879804161, -92.9260669123227, -12.8877098522159, 11.9254708708532, 
    70.7248759223067, 69.6138198488274, 69.9365169623486, 46.7681351237052, 
    70.0025907206241, 35.8881327687888, -38.609897563662, 41.8579210131353, 
    31.8047821558349, 14.3632082437022, -26.0012795354926, 19.6093813036258, 
    -48.2593835155513, -33.7115627334636, 59.5241320363494, 80.0247120501998, 
    47.9091484347195, 13.8505236803262,
  83.4419341946317, 12.8192376110014, 32.947292008976, -27.8832997998002, 
    -38.0301524387166, 19.8941913468795, 17.302227585631, 72.0245781451906, 
    22.7096367691334, -0.873197633840973, 19.8380373650435, 
    -55.5414273312137, 70.1742677244438, 2.59865913227215, 9.43834717446019, 
    43.6080148645748, -12.480880009814, -28.9842184122003, 29.4361331240987, 
    7.41388694424071, -18.1849365343824, -1.83047080537298, 7.93982483374742, 
    82.6404176322941, -52.4781579601784, -42.7331377839908, 63.0278901472804, 
    45.9326260751171, -5.69807685234739, -70.8280220949158, 46.6399771718807, 
    -74.1636869068064, -42.1969880893501, 69.4016543439787, 15.5049415054865, 
    -5.79617610792511, 105.090482846013, 39.4677305827395, 80.2871365587365, 
    -44.2629594389538,
  117.341268761216, 58.1676996078712, -60.5841834201846, 6.50609690734226, 
    20.3488061312134, -98.2405413283671, 22.2774583859915, -77.3346608459928, 
    -21.6125281250999, -1.03315497253812, 7.98627648177921, 45.1574755979337, 
    -87.3115184806865, -32.9360589217216, 39.9958111331848, 
    -9.00129984322206, -8.45800420098179, -23.8860869367058, 
    -40.1215178129024, 25.1110779903616, 64.8165292520738, -42.6083038324299, 
    18.4011486504478, 29.6819873051123, 13.7291166704042, 39.8583907586296, 
    123.218083242139, 4.03575653892858, -16.2973600230004, -5.19232231622975, 
    40.6842342551607, 22.9790409541912, -13.7857612192484, -7.67070710510564, 
    -16.8060594675605, 34.8244879201053, -14.7681282805717, 
    -52.6107368655511, -99.8703479924392, -26.3143115588315,
  93.7525778318715, 75.3840894262199, 77.7719903681967, 27.9654740974461, 
    -6.36377463281334, 25.4764833536284, -37.1327665095997, 68.8386261655254, 
    -14.5277852537353, 23.866212961031, -35.1534942319111, -36.3682962488329, 
    -44.1281009778344, 73.0997833991458, 43.161021333244, -29.8634814864546, 
    2.25274212954386, -43.3086276264331, 104.06919544201, -15.9066816246492, 
    18.1506396362243, -69.7981878287873, 84.0719515190498, -81.7226959180528, 
    -36.5105762883477, 18.3331842944347, 58.6421336825319, 14.5100059988066, 
    1.20451208903118, 22.0329507194702, 109.938748125656, -62.2595514828079, 
    -76.1876049492596, 65.3104341650732, 102.578141989021, -64.9348796948119, 
    108.382823699958, -8.19332710487724, -27.5789562431981, -72.7897820529429,
  78.6537459612272, 44.747105188565, 33.1768326853481, 38.5199862187549, 
    -36.975141423143, 54.470411562419, 97.5941169938529, 4.17323303165537, 
    22.0607295893333, 47.384412947766, 0.253048218069951, -8.22687788179171, 
    153.058568519049, 12.617497040344, 32.8510755006545, 31.5445750658238, 
    23.2108862292802, -1.02485668784104, -52.5779175231115, 53.8242433827816, 
    25.2238249091142, 82.2028390069847, -8.24656060551897, -71.4604694732913, 
    -55.5861671878438, -4.2809036151268, -1.25370125863669, 51.0659739165691, 
    -32.1204504524761, 2.54025339744572, -32.6425314566878, 74.5045327945958, 
    48.9712337696553, 22.6047832595999, 75.0912565049164, 27.7694597863359, 
    -24.9322706777578, -39.5480219392401, -25.7347891980737, -105.48187101491,
  -10.570137028959, 62.2332842042102, 19.4458773521105, -17.6255007724019, 
    -14.500030773748, -78.3212880201339, 61.2790702484512, -7.65865963184134, 
    -28.377267462974, 42.5252311859726, 25.9456039684848, -20.4379410025373, 
    -96.7026838866705, -17.7448936519561, -26.0220146915989, 
    7.45959322575232, -20.6795358330234, -42.7890046109237, -20.112886401464, 
    38.5003273269002, -52.8517340805329, 35.3851599785638, -49.8760210640117, 
    4.79120185160626, 70.5600719645423, -22.006819470257, 27.1749948673559, 
    -44.8821601653676, -82.2014021480446, -3.18510254559426, 
    -69.3416447311879, -48.9295291797148, -30.3681211550476, 
    22.0598519950148, -3.14940051201646, 0.471262939617314, 13.3351672314312, 
    63.122728471316, 31.914157409782, -63.0589469854782,
  89.663065715384, 5.78023592452037, -12.8109945098981, 38.9137612355278, 
    80.2401099235628, 50.1361016559534, 15.2492100449623, -36.6433828473102, 
    5.23139720191958, 54.8132290669947, -69.8264836928851, -40.0051523228326, 
    32.2015718362087, 66.4521115169079, -2.15119479160937, 33.765682129213, 
    -87.8930463743659, -68.1196200133597, -60.8951377771658, 
    -5.92502367354642, 29.7106890338507, -54.106630110195, 23.4557695243854, 
    18.8113452740856, -18.1279273804572, 75.1699151001794, -17.1621429194314, 
    -95.9490872571765, -59.924426771044, 53.2735481119384, -42.3947241087524, 
    42.8911364907831, -50.3163651965153, 12.1182902670008, 60.0702304141961, 
    19.7636817716036, 49.8483862614585, -10.0200658818188, -43.3858577362027, 
    -14.5326197186719,
  73.1237434742565, 9.58079737104954, -15.5299179645413, 31.1940386783351, 
    -15.1444658231904, -7.28641754604888, -22.9473950700033, 
    43.4587842572026, -40.1940150829061, -73.4018170314844, 
    -25.2988991341989, 100.014927400626, 109.246202906243, 60.3585778031473, 
    48.1125772049453, -23.54696874446, 10.559410771856, 68.4441570670308, 
    145.299263953664, 60.1670324588049, 24.2389091895995, -32.4480194554765, 
    24.051817366963, -18.782707074988, -21.994934808201, -14.4823507685697, 
    9.62885314058108, -40.8749152656887, -3.58787694751252, 4.86679718981207, 
    49.2684014433695, -79.714749980023, -15.6745958266634, 81.9373832458752, 
    64.7724561236352, 59.3837464337309, -13.5234965173299, 45.3217186538554, 
    -43.3931197785203, 40.596019259843,
  28.3313152613037, -81.8751577101383, -48.0842652923419, -13.6991118926227, 
    12.4944237201066, 80.2812951975671, -63.1305546150262, -14.6858552044781, 
    -21.3638446489365, 25.8045727944374, -54.9378882010474, 
    -30.9168190261907, 30.0906204407961, 33.0611203735938, -57.3728530977324, 
    -54.6975360082489, 39.9981702849913, 66.7267572034218, -15.2515209306005, 
    -5.56256667190113, 59.042062728114, 26.4614713733512, 34.1310819140653, 
    -52.1708826185598, 87.7569895211755, 31.1069022081631, -3.59785523706255, 
    -134.499764954357, -4.48651614480122, 30.3158646586285, 11.0350949468734, 
    7.34987584492133, -55.7985953508243, -87.8783862133843, 
    -36.3182664231892, 29.5492087935724, 64.553751457972, 135.366084565882, 
    -34.0130858069595, 33.506254087099,
  129.225551375186, 8.36807670177898, -5.19329768580718, -7.47863337527997, 
    -40.9767018767749, -20.3418992799382, 38.8845596295178, 
    -21.4595010135219, -34.7445637822394, -37.1900452777241, 
    24.1954977366415, -31.6899771655804, 79.8557275850009, 2.88714214167531, 
    -21.2733236116642, 0.00224001206519761, 5.36103861265471, 
    -52.0644007848065, 4.99476888118875, 26.5733743472957, -14.858217780206, 
    -52.5080264829514, -18.3609703110941, -53.0905501183217, 
    -50.7397808134813, -89.3796129498373, 30.2591400460755, -35.779792301653, 
    11.8056317716386, 69.3280411759789, -80.3660975714047, -30.00113773456, 
    -117.703882615006, 57.2585823849903, -91.3526649956536, 114.624006042245, 
    88.0634325182214, 9.11185779837236, -46.006382294454, -6.94345167687287,
  107.53308751982, -3.79830251517696, -62.0422115878187, 3.72358669039883, 
    53.9278374236582, -3.10572257640848, 2.68115954127726, 111.747334757874, 
    -57.5529018503721, -60.5667279034612, 37.4448628869582, 
    -12.7042022148935, -50.3728626529654, -4.72165588758351, 
    72.5218660133638, -28.0616865580825, 48.8031502542679, -48.1467068359209, 
    1.51736802017111, 111.808593769614, 35.705302256275, 128.040207502587, 
    -61.8099837435351, -66.8062707679906, -81.0332594729065, 
    57.3615492923337, -71.9766387320204, -82.2155683761477, 109.577057241492, 
    47.0999959670414, 10.5404596290201, 101.137134179344, 60.9830444596401, 
    55.3285371473574, -40.0969379315468, -91.149959820054, 32.0209777518512, 
    4.96600419096691, 11.7546956067177, -36.6366946102467,
  91.7593153999689, -19.1229841213491, 10.3861994001968, 56.892169283227, 
    -2.87731730829394, -8.26684172500148, -4.82273365377971, 
    -78.6148222050284, -12.2342149320816, 59.189918829961, -7.00003684497495, 
    17.1567179761521, 47.5943961735119, 2.39991593274146, -49.7658894982023, 
    -6.4797462312957, 11.2941531641998, -43.9728514362873, 97.6064464377662, 
    13.2838449751046, 57.7595140954096, 37.2672062618294, 22.0520006273972, 
    -102.288872122168, -11.3816208258543, 11.7558973031022, 35.6025684845373, 
    118.272196635883, -49.199727392318, 42.4361565511346, -19.9048896350969, 
    -7.23738419806019, 55.7274421860919, 7.68669758859856, -81.5439514948992, 
    54.127836117543, 1.5506429321724, -16.2263020260888, -16.8461144104322, 
    25.5712717188385,
  97.2878465029408, 38.0147451933253, 10.31540193886, -130.996050464948, 
    -41.3835021646236, -44.4904759767809, -96.8510976103085, 
    -29.1577731831858, -55.1980038215334, 23.5653894744667, 41.2658045156176, 
    -71.7902934909777, 72.8647849040141, -89.7572012208706, -26.320146359999, 
    -13.8493082000345, 24.8439380124302, -61.0496551896847, 
    -8.01632683183056, -13.3405774994098, -7.55195206536097, 
    15.8618562994111, 34.3155776630782, 94.9675783879264, 116.839248190667, 
    -37.1301212317087, -40.4422123948029, -43.1294042099968, 
    3.47513110900794, 47.0227871598336, 149.755931502636, 5.90341353392892, 
    19.8040053197049, 20.2746557072616, 45.6796287907417, -29.9956445339101, 
    26.9732278239815, 12.7828563162544, 44.4072654760365, -48.5913057339193,
  89.9098114674495, 76.6172705344624, 50.854262777026, 20.5981176170615, 
    96.8637395968501, 52.926373477028, 53.5056545042916, -17.3468548986348, 
    32.5272813085291, 57.3886538479356, -60.2954785396127, 1.4360946280672, 
    -20.1494731188238, -11.9129130134648, 24.4766733413093, 
    -50.9498657679859, 22.7955908748031, -8.87642617437677, 
    -12.3728003032633, 45.1190183620936, 49.3357430617962, 12.431609919783, 
    46.2293033469956, 27.2063774255119, -60.7326123840563, 8.2823107772816, 
    30.165065143759, 34.1413703769123, -51.0933089796492, -17.4762566986692, 
    -46.1667919316227, -14.6702219620224, -16.32557432038, -22.9208017285369, 
    95.050042749405, -100.243824426556, -81.4914496186455, 95.739359867333, 
    -19.3093619905319, 52.2923829514361,
  143.885436728213, -23.9567566593777, 14.2674828460505, 3.93675190091194, 
    -9.17934585919814, -19.6620539600532, -30.7249122290371, 
    -19.7777889332402, -46.9862411973071, 25.8977339880243, 
    -76.1302043451292, 39.9808196013502, 98.4375469181828, 26.8014061920283, 
    21.4714205014495, -72.0842987724973, -29.3092923361856, 130.328477193222, 
    -13.5324435184317, -43.7473962508018, 7.39991513633827, 
    -29.9211273745402, -17.0369755001618, 94.6865805090321, 34.2329749946136, 
    -52.8537739417462, 31.9227858511002, 73.6879174379034, -22.3363909538607, 
    -5.63595995269285, 14.0703601646807, 66.387752510756, -11.0147239184954, 
    60.5945374722876, -53.35612241634, 18.5509990724916, 59.2329610182459, 
    -28.4268906984519, -31.3679900838697, -31.4704281216366,
  136.576797325752, 1.55867883453997, 60.5603290439305, 21.5056262036341, 
    102.367165218632, -27.6518486979916, 2.59025923679764, -43.4267046790777, 
    15.7100608776674, 28.6721278946545, -21.0365014179434, -55.9083298248001, 
    -43.4423237973456, 11.5879711624088, -31.2156900474727, 
    -6.34818219860963, -15.0250950383578, -71.894681021406, 
    -44.9640125519749, -46.830193408059, -67.1060988695954, 12.0438222981097, 
    5.07259467216129, -35.8860734275581, 50.3668528722759, 26.5165854402449, 
    -83.2995283209444, -63.7317530291577, -31.5069097547308, 
    -2.37676714320359, -61.9059871043622, -27.9303896517691, 
    -40.5666278447201, 34.506124134298, 7.35220741568416, -41.8276603436882, 
    82.3557122893165, -28.9128984901185, -1.12342805580463, 11.0678099298408,
  94.4508287287249, -36.9896181419132, -74.5154118253226, -18.3742111717292, 
    -39.930871091158, 46.4664075505778, 100.185357855491, -11.5622807200094, 
    20.8645071769074, -96.979653355903, 70.1193039147434, 49.0270767787055, 
    23.6726736986393, 7.43768958941726, -15.0036650719727, -30.4672735782854, 
    44.588919730441, -37.2873064665588, 15.8357190605746, 83.4576258764181, 
    1.29139268154332, 116.85622335156, 48.4376779427087, -59.8354668973695, 
    -18.4275898748341, -45.578449035386, 0.798685412630113, 77.7066554359879, 
    -38.143127509789, 3.6448212858992, -20.8977391261068, 7.52847006463209, 
    -3.23604699290054, -38.3084594931564, 53.5348635856705, 
    -27.8462306207599, 61.8336496905448, -36.8418060581573, 100.199787088795, 
    -6.58947290562223,
  132.383558765994, -32.332981623065, -78.7847448136141, 31.0151413751677, 
    -60.4547432999892, 82.6554978855789, -1.30696000227047, -45.548960472381, 
    -52.6909566186774, -8.69246607038319, 108.797315028829, -74.285779635333, 
    -29.9837269475888, -70.812976569092, -103.788352332795, 
    -38.2767700973077, -71.2335171779884, -6.56316757376533, 
    30.0508891102866, -70.664028906868, -11.1946089579593, 24.9262241318108, 
    -3.43304870706775, 24.860918833714, 43.2011689642887, -28.6194047745376, 
    115.977715011568, -46.3422907610032, -6.56263974240288, 
    -47.7663304131896, -31.3898340379669, 106.309801226547, 
    -73.4680925615535, 8.31833499862144, -43.178450031423, 6.0468128549535, 
    47.4502504106133, -9.40483092686852, -87.0757653293854, 114.757771887042,
  73.8438131070587, -48.0470747568972, 85.0795956480746, 56.9782450299084, 
    51.0102197575882, 46.3656000016837, -40.4310505850471, -4.33457054019362, 
    44.2602416138128, -17.9659265519509, 42.4303728957474, 89.9765296103004, 
    4.07827070314929, 94.1501193108095, 131.786561282263, -22.1817380582871, 
    66.5118841453394, 94.7128173606572, 11.5642572446975, 12.3537531157678, 
    96.8518945837591, -4.89161397691609, -42.7644218395462, 
    -30.6281091317426, -74.8564839841676, 23.7936340841231, 94.5898934197274, 
    39.0090679982165, -75.7560155388912, 6.32743062514255, 63.3720722919196, 
    -85.1390017967366, -2.26883500868958, -49.6803329364937, 
    26.8766653470773, -51.9638102478855, -26.3262337049599, 63.2115559642422, 
    -40.5531816711467, -3.86671356472075,
  108.636650460641, 21.4034000180035, 77.6967559440856, 39.8948455604526, 
    -101.10056633163, 45.5544799786605, 30.0742640214759, -94.8888745561271, 
    -52.5472155369882, -117.404899130813, 24.8463649924698, 
    0.876815141227105, 0.989636256488464, 25.1553095669049, 
    -6.21472938844509, 41.309159058899, 14.7565160602713, 155.774442554598, 
    40.7930807018808, -58.6306744037599, -51.818756655741, 1.73118510075954, 
    78.745929751182, 138.291844296884, 12.3463634880543, 5.62641187945859, 
    11.8298942195532, -6.75985323381391, -1.76537658752858, 8.91554012539723, 
    11.7227287076118, 85.9368279891876, 30.1412902990382, 11.2222761965108, 
    -62.7519497959086, 61.1491216205907, 33.7292209328219, -7.23244192636517, 
    -26.4125566723179, 24.9195602556983,
  123.831311583312, 55.9359351415764, 84.1118069407671, -22.07771767369, 
    -34.1750034474456, 78.88323240335, -37.0633006074475, 91.6478522297815, 
    -4.10589260310348, -61.1301324082496, 55.0472853851057, 84.052138377743, 
    -112.214399056155, 31.9461265854845, 26.5634485305219, -15.4229071661975, 
    -70.9908396728656, -13.9963206916552, -6.48220753891256, 
    -57.5243429985599, 32.5568830571444, -43.6677459103103, 45.6371185739597, 
    16.4311081309837, 34.3991420125575, -21.1650708632471, 6.60773192287587, 
    -26.9889369546482, -29.9462264543728, 10.0685389727525, 
    -82.1059892458214, -47.209152765524, 23.7113146810634, -33.2957121645292, 
    -5.5653518535795, 47.3027593568054, 15.4231250762216, 26.958352976692, 
    1.79364493413396, 27.9742894243203,
  43.8024576616104, 16.1155089842768, 45.3620884634113, -30.2953776651429, 
    -36.0913998846992, -72.4415222041885, -11.7494126751733, 
    -16.2595219816765, -40.9558457812582, 38.7825779772461, 
    -112.058857633793, 110.75136091159, 79.0085186989873, 13.1959969358864, 
    -140.143838362531, 6.39249303923494, -5.6114584174778, -67.2059107945611, 
    -36.597700041652, -19.7298183188973, -33.2828853141591, 72.5336729017605, 
    79.8989907258899, -33.6948915554433, 3.18256175132931, -81.8446118766609, 
    135.39110642484, -1.52424957313134, -41.0980061338567, 15.5664763060347, 
    -59.0590671211055, 6.53319727740088, 39.9338978484872, 63.5036270591163, 
    -54.0179316873784, -56.3400051809107, 7.538923129271, 91.627431560174, 
    -120.598250720536, -22.1756045748714,
  143.056360703103, 41.7626935432879, 108.501333948762, 5.55600823265403, 
    19.9861805662339, -2.17887124716031, 56.7959534197491, 11.687481436309, 
    -214.48036505689, 51.1527752393715, -13.1135011928019, 88.1863784854201, 
    55.2562468445509, 40.7075029304013, 47.8823375655085, 17.5357373986827, 
    -61.4921393234536, -62.5979123661745, -0.609122866285409, 
    -47.5892244829722, 1.51249853159921, -65.4962997676752, 
    -28.7751210886468, 42.0718386459853, 34.1821028872176, 60.9005997149997, 
    108.556548153581, 39.651654045301, 26.4641775145276, 65.6987120327273, 
    76.356882332664, -67.2956563055141, 104.246861656209, -96.264914248953, 
    36.3526009594197, 41.2254514699776, -23.2711409839622, 43.9338921094983, 
    13.6328675700276, 40.9282995202757,
  100.436635192605, -39.3001260591891, -7.28411021104527, 20.7497048300138, 
    8.16757302992911, -38.5776700600719, -40.6189804111571, 136.812640120604, 
    -62.4401893535686, 28.9990034014958, 46.3605261427681, -41.0762220755923, 
    7.79765840428851, -21.448260889828, -74.09243316289, -67.2904270603761, 
    -54.0578604554775, -50.3391641001174, -50.4346702195558, 
    31.0264341064884, 10.7781213289572, 29.2632438381052, -15.37168530127, 
    15.4142772490342, 64.8467241437064, 25.3931067334742, -71.3992514914541, 
    -108.479735231398, -97.0774577575141, 71.6567445709777, 25.1942893055642, 
    -99.6675301476969, 59.4139153908301, 11.8300775518014, 3.62719620199087, 
    20.2906467736697, 9.36005496752605, 12.0388062546388, -52.5789366174702, 
    -42.3280898294544,
  62.7211610126714, -1.21608551723786, -15.8844840286693, -90.2724154789737, 
    100.128177066948, -51.0053727545786, 18.1172759568858, -24.5818573949896, 
    -30.9069982962065, -19.3946260642463, 10.7369458354373, 79.088191272123, 
    16.0759147873415, -35.7478692208399, -56.2034902149983, 
    -4.90319728876845, -8.20639497024374, -50.8411781577892, 
    -4.56359083278417, -46.770315861489, 62.771276742212, 96.7941078016511, 
    -59.7919481545649, 6.64400609605118, 92.9233899226623, -11.339678588469, 
    -27.4914416673587, 64.0479715281205, -32.9916016655105, 8.7530807206763, 
    13.9877455573684, 53.3249111988788, -5.52889877293979, 39.0202624474549, 
    -64.7261081007165, 36.2703348626002, -10.767972868249, 49.3164287004734, 
    -57.7594796783072, 10.0775241387304,
  119.161460118091, -81.0464669433908, 38.8019260934782, 58.8998457871467, 
    42.8916060401154, 104.203726943062, -17.263101766404, -88.933819391986, 
    -47.7135244359215, 19.3092924903722, -34.5570399593971, 9.20220419299649, 
    82.5041115019902, -6.02503718498006, 30.625515593188, 30.6085316908213, 
    -20.3972516307024, -2.38506835636571, 39.1783399156012, 
    -12.7321582703155, -63.0661932798169, -5.46504755699289, 
    -55.3416918737173, 12.1571737504079, -34.9453225580686, 
    -26.4603394047084, -0.756310341079615, 3.4204153146828, 46.2474751705467, 
    83.2540673456699, 104.41188410428, -13.0485821104666, 44.7532459895909, 
    -1.46124350522094, -13.8861833426369, -20.2075890819419, 
    -47.9744339868901, -76.8729658799403, -15.0637469116615, 23.7121820861809,
  139.984179464291, 77.2689372086907, 33.1527312346599, 1.18687071165455, 
    78.4871325765673, -107.139575499817, -106.020923524977, 
    -40.7669096108947, -49.1842249922427, 3.73648383032173, 42.0908460082749, 
    19.0664404300949, 42.628564621577, -37.7795922805845, 84.260424778355, 
    -80.7592355644838, -21.9255710026694, -2.58144913243031, 
    85.9404215257159, -32.5866957635276, 1.08531963664384, -4.36256167659345, 
    26.9587282309665, 40.3919698664098, -43.8204070648994, 59.4983917132156, 
    3.22335819840241, 25.4531670895536, 62.9290226268267, -31.023421529865, 
    31.3280122353147, 24.6350330509061, 21.102924802202, -68.7763577104246, 
    31.7570438973592, -36.2794691982221, 21.5180698056161, 39.7261892596027, 
    -37.1174789124846, -16.2097639329527,
  142.224433005994, -34.7154106656952, 1.085895699096, 87.316992717236, 
    -62.5519804431161, -28.9794473841162, 41.7823585376166, -24.118260095588, 
    65.4629201971573, -67.5262964161962, -57.0737018427116, 25.4718243251753, 
    2.62991736688329, -5.98400086988745, -77.4148625515317, -152.67648892581, 
    19.7756497866953, 28.8282138606741, -26.8902035154227, -18.9144482509372, 
    -18.8061692057143, -35.55066216157, 4.18798378643675, -91.3671390881375, 
    -0.543569129672016, 3.39425580843941, -1.10046861534322, 
    38.0995994905164, 8.74449282495462, -39.872574693312, -64.0114018672525, 
    -16.5374908023249, -49.865126735886, 12.1237837010679, -30.4193315947401, 
    -31.4653926757365, 20.4911638373033, 32.4960376167011, -47.8372202652327, 
    28.4197085696719,
  177.542377855523, 2.14071854957114, 32.9677508027906, -17.8733338078774, 
    25.2099022641349, -54.5926125358989, 14.5717753260188, -14.4990014337256, 
    -26.2025687490598, -15.9959423908836, 5.90258227273848, -45.389741523395, 
    17.1263065836722, -8.55213851360028, -12.8896500061756, 9.54607415800682, 
    -64.6268216177814, 53.1960615389952, -47.8038153056711, 41.2061656467741, 
    18.2201048812389, 23.5266377287494, -11.5536671653406, -8.63429771573098, 
    35.918093787735, 68.8216286026009, 37.9307236419539, -24.2695695163757, 
    21.3587644271641, -59.1642167399252, 86.1007747705341, -53.4388668105642, 
    -6.02753163099797, 128.012972035943, 37.0611745928819, 49.9099713754881, 
    -104.195285224993, -70.5736872358281, -38.5314950546117, 75.7144928112149,
  96.1353438151707, 10.881269324296, -85.0746739858665, 35.0711386140879, 
    -28.1726247547871, -0.75576445886017, 18.8075655417094, 11.9793930170004, 
    -11.487387508082, -43.3801729265621, -69.1688661610467, 3.94053838001589, 
    102.628611069256, -18.283869855649, 73.6545789835365, 27.4006445616419, 
    52.5138004181375, 21.3867318527695, -15.6881360859384, 12.1891763187408, 
    -40.5346910257147, 84.5320847224389, -11.478900057445, 100.532538548209, 
    -12.0591397711084, -14.2586245179095, -76.8011479202886, 
    -67.0593831739722, 33.0476732510506, 17.4166664510208, -40.0134831397678, 
    -16.7623665725252, -113.924085706463, 89.720910037824, 4.98804429162574, 
    23.9709522362781, 37.4199471335616, 11.2263799409359, -10.5150358907257, 
    26.0907865334714,
  224.874824737533, 117.114776387573, 12.4921282872316, 7.15004388077862, 
    20.5339165035819, -22.7347848157449, 17.8536316051751, 36.0061916742813, 
    -0.165750604727533, -13.1237007421276, -41.3529221471804, 
    -2.12513589668118, -48.7326885841406, 54.1424267809303, 32.3242433491539, 
    8.98462910654369, 37.2062192007577, -20.1653154539541, 14.2527213084806, 
    -34.8573237013675, -72.8080464354784, -44.7504631693117, 
    -97.7800752765345, 35.5134734028696, 81.450190036039, -1.21081308262836, 
    -39.971827770634, 24.215703933173, 12.7772846530878, -6.38984818323976, 
    -40.3494071416455, 54.4192125045037, 23.0840444878246, -15.8123935799228, 
    71.0926659312979, 52.1631159419858, -36.8516363893249, -93.6691487897995, 
    77.4765306585459, -18.7035009189386,
  90.1652961464957, -15.045038250904, 26.5314517393484, -5.41585785941517, 
    35.7766775146275, 31.9490973653185, -71.885737662474, 17.1733544423999, 
    1.92381256996499, -1.86149001850629, 66.5959695849872, -1.86345556251358, 
    -41.0649974652271, 22.8919013334642, 1.10195696844952, -9.49159912316267, 
    -90.9923025426792, -9.51589159217834, 29.7622065018935, 36.1647534585807, 
    -4.05138131989181, -40.6987482356962, 39.1603563650906, 28.9070663549448, 
    8.26336453318478, -20.9746572578183, 34.8414005442677, -5.28850867680115, 
    68.5152952495663, 24.8293600128783, 12.7763884040104, 5.96182655687794, 
    -62.9100735001791, -87.7838437200495, 42.4345156547699, 
    -52.1693446234333, 61.8078339433552, -39.2871825545269, 66.7145951443491, 
    103.018178343819,
  16.9114766063556, 16.9279882444826, -56.1348337160195, -86.3982476985994, 
    45.9620611801341, 19.8958707413066, 69.0594884767051, 61.2771482901596, 
    51.026600897928, -53.9741301788574, 96.3612660297935, 6.54620283346663, 
    33.8579727727505, 9.81462732891151, 12.3693062677693, -47.2053787609714, 
    83.1690849717893, 28.6718777782262, -66.292121625551, 17.2972828391465, 
    20.1936913943621, 60.5215107281311, -18.4268590776672, -56.503552721349, 
    -73.3171693752992, -80.5240209040222, -41.5684178571484, 
    -125.339134519502, -32.7669642043195, 58.0000845971454, 29.0015883047268, 
    66.1860791786065, 43.6323103553827, 4.81787084193119, -64.0068264544069, 
    90.0155132706609, 1.65644017786526, 3.03035872432106, 40.2717120860964, 
    25.9361802146513,
  24.5207401369313, 48.5867990916099, 38.3947583779559, 24.1015799107561, 
    13.2915558813444, 42.8270552111307, 63.3821708188304, -19.4190454630639, 
    -71.2477600578139, 18.8910484814175, -60.178806301607, 35.8129096017297, 
    -65.5766588414768, -92.7999235087899, 37.2097350405304, 
    -18.4451752307834, -2.49054732953098, 0.438175481513156, 
    19.7178699267834, 84.4138700058397, -25.7446099335086, 43.6958188159625, 
    55.5352929829856, -51.8951847946521, 19.2316827627895, 33.4687172513696, 
    2.80823540864655, -72.4944791875707, 36.085517099328, -73.8648173147041, 
    73.6736848725131, -50.6687559331071, -2.11474806742685, 74.92701074929, 
    15.7101777604594, 26.9058615692527, 18.7499518464291, 15.52053295233, 
    -26.8687626036401, 25.3128446895972,
  132.419765335543, -43.3686638626918, 60.3435554822251, -11.0838444112653, 
    36.4475167744647, 32.012316680633, 18.3402919923829, -62.3820572028814, 
    -81.4070512403515, -77.857795858616, -20.3953113106716, 
    -59.9329954462857, 3.69687909756875, -5.48998497735334, 44.039359442915, 
    77.4468104032361, -81.9041002922656, 37.0733067498916, -44.2452179786932, 
    21.2740442791702, 77.9679107421268, -71.2252549377159, 17.5731684545313, 
    53.4822133858167, 19.4842763646963, 113.160716067952, -66.20295800839, 
    45.8103136660662, -7.02209947442169, -72.2228608075554, 43.548475765401, 
    -0.0863144210642136, -67.0137875979444, 107.341782339179, 
    -11.2758197411418, -24.5372971472191, -51.1401133939005, 
    -13.5773865450659, 58.0697400392906, 16.5069603346171,
  128.855669572704, -10.5567241809605, -1.01953125801595, 42.4674721789961, 
    35.2243894655491, 27.0897653664082, 13.6551943987383, -57.6145230392089, 
    -47.0894256709309, 29.4068154312759, 27.4793901348777, -29.2355557936533, 
    -47.8370019157456, -65.0668243705408, 50.9988238555354, 17.9441974348137, 
    -16.3274114561327, -35.3805829294535, 0.0189207175193777, 
    -6.44445889125014, 36.616282765755, -53.8959182738554, 49.5415673956234, 
    23.9244935040578, -16.5844855622026, 1.66906516816867, -38.7510982938555, 
    53.26477139268, 20.9017707388471, 13.0187526595734, -5.97640487210627, 
    -4.82275810179447, -33.5434824574365, 100.766672683435, 74.2554907054194, 
    -41.4975762441128, 58.4564639239961, 65.5091274383946, 46.2422584557214, 
    -36.8684442206713,
  146.758177416116, 47.9350810504338, -7.66730390890906, -14.0216227426476, 
    -31.3793706724785, -98.5552506948366, -10.8766992209046, 
    -27.9403993651407, -31.7392655617256, -89.0180789213517, 
    -6.54913696715611, 100.478694366197, -45.4080765525782, 
    -46.4341352613831, -82.6336853049886, 20.9543015292153, 114.603157222837, 
    -78.746865495764, 37.2706284258829, 43.6572848837776, -26.7673983252028, 
    -37.5113642100205, 90.6880737739128, -99.4189813717228, 
    -10.6515432837607, 15.2735834942749, -31.5937314495211, 
    -46.3525554240666, -0.77993434620172, -8.39202460297164, 
    78.0513943215569, -4.83898292938679, 50.7912663258143, -43.9290925366213, 
    -19.7454605235804, -61.7576283775453, 3.79925935491965, 1.99363014516768, 
    1.96341398782758, -38.4624637581321,
  103.1438717241, -90.8359923342933, -35.805320933045, -15.648783298216, 
    20.3906059296824, -17.3810182814732, -56.9190653994995, 
    0.241933507755392, -20.0990484782042, -30.1583592543345, 
    -39.4883377865023, 7.50163631137013, -49.2438473166611, 
    -5.77427551242768, -27.5641304677424, 27.1803504414323, 110.929297928414, 
    35.2313170925569, -15.6577622788012, 52.3157935136833, -37.5276775253567, 
    73.4038822363623, 10.4202593092634, 62.1984463113654, -67.4245353477938, 
    1.24606605577671, -32.9801890831883, 24.1953671328897, 9.27972748930368, 
    -52.3613098930189, 7.70480331200191, -10.4781391133855, 43.7511088621835, 
    8.92113032408897, -19.0015329610996, -19.0799877762085, -54.186305952972, 
    -48.3315527262056, 26.3339968748511, 4.14356848936888,
  66.9781938932997, 33.4464306766185, -93.3704015673846, -9.74916537706952, 
    -57.9708560058556, 18.7514276457301, -11.4986937434666, 22.9980674982227, 
    87.5142458324863, 19.9041167708245, 14.5819380215534, -11.4399374859331, 
    4.39787498727839, -110.629898276785, -31.204704606485, -7.19061604684047, 
    12.5778809361505, -22.4014398007617, 39.2026615080661, -26.8467646756954, 
    7.18365180292831, 27.483218204458, 29.4013705937393, 5.15998113936346, 
    77.2655630120965, -25.7273650892319, -83.0253029056644, 25.2284367282355, 
    27.7449613117576, -53.3962965438387, -46.649056391881, 33.0480474211255, 
    11.4121835436789, -68.7957915865151, 50.6482614794969, -3.27618793581882, 
    -16.9122397355602, -21.9937458301808, -69.8741646095177, -26.221836424627 ;

 state_variable_mean =
  1.91656620796571, 3.66785779883771, 2.80447246024572, 2.14256780448976, 
    1.83070186080589, 1.18898746266785, 1.88930720316563, 2.86504596157058, 
    2.62091679584613, 2.78499701413629, 0.613585153421966, 2.30097322975582, 
    2.87464026811012, 3.43783106692137, 2.84620107296898, 2.25410755916963, 
    3.05385563819217, 1.65269884735824, 2.14933974382213, 2.19788171818385, 
    3.43343596080859, 2.98147433096104, 1.54248829020696, 1.75218747195477, 
    3.76172429071222, 3.09968534885687, 1.0943805589739, 2.01683485399969, 
    2.75281912038066, 2.87200260848951, 3.10324839686578, 2.30507051298501, 
    2.79993614208648, 2.49850566474607, 1.76329992719109, 2.65037691532444, 
    3.00820397461436, 2.19961686281177, 2.42443072161339, 1.63959947530192 ;

 tracer_concentration_mean =
  9.20699946725049, 5.52428721186081, 6.56164065076612, 6.37290513830332, 
    5.8303813700075, 6.19093794597121, 6.05547802297737, 5.96381919681991, 
    5.24624368960605, 4.41892921467131, 5.2466911692408, 5.36263736740687, 
    4.99934342046685, 5.43422936548071, 4.77890511873222, 4.68587169661648, 
    4.62345339315521, 2.93994099656443, 3.89074160734733, 3.71676808330054, 
    3.2615455773603, 3.83048309475909, 3.7557994082178, 4.02869317741781, 
    4.20135249251821, 4.76596345804256, 4.82274232735643, 4.18232297894917, 
    4.04212418937996, 4.55114895779149, 4.74361719195326, 4.6440695461851, 
    3.72385796017496, 4.14367531642239, 4.28314215814055, 3.63543902126022, 
    4.11056500909645, 4.33641071692418, 2.36472141760282, 3.96614222884049 ;

 source_mean =
  103.186573147602, 7.90073070783628, 6.71471350792824, 7.04236688374077, 
    6.72865950302913, 2.42277169693692, 4.21819189076818, -4.11747360613053, 
    -21.4399428960998, -7.6260936302757, -1.73485117247503, 7.48992299555976, 
    7.07966970696598, -0.244660071210813, 0.392842889476322, 
    -7.58263120698046, -4.07900797854915, -8.03862124215612, 
    4.78618288478314, 4.03338762610633, 4.39377652919019, 8.03200597971819, 
    11.8126231757514, 4.37337183650044, 7.3205501247594, 1.40365630843318, 
    6.55927525132577, -6.12890942517463, -6.56275595186466, 4.46837932544796, 
    10.4523095301459, 0.941867406263773, -5.99684158633523, 14.1933595994827, 
    4.1021520225219, -2.04172456470127, 17.493755531805, 8.6749379413066, 
    -8.48480661699252, 0.51690928017398 ;

 state_variable_sd =
  3.35685155081193, 3.81935520117529, 3.85394478448017, 3.79661891868788, 
    3.54049723335225, 3.58926402508787, 3.07939976980902, 3.54022415908232, 
    3.42321134246925, 4.46289136514446, 3.28782842044213, 3.91758834144164, 
    2.95327671712543, 3.63961862487362, 3.25013223244737, 4.00684857495891, 
    3.49787310194981, 3.52901346088387, 3.78282548884337, 3.37287866929827, 
    3.59752825606075, 3.59787002942786, 3.64803382151679, 3.44268967649971, 
    3.88014524928764, 3.93649264640168, 3.18086608596702, 3.38417153206127, 
    3.65922615477097, 3.36812680307808, 3.52872084870505, 3.95213443381477, 
    4.05777840735479, 3.7218498155839, 3.47055709676415, 3.33738488779088, 
    3.42965584589997, 3.15748185858822, 3.79862429103676, 3.68703675423544 ;

 tracer_concentration_sd =
  9.20496755632266, 9.26285869501813, 9.42692546017446, 9.19947788724431, 
    8.96585106925265, 9.78896311165326, 9.65139859970703, 8.67155409136191, 
    8.3921961465199, 9.69342013379207, 9.16724390210143, 9.98303186751154, 
    10.0865414811826, 10.2679199321581, 11.1272265525434, 9.73595095321427, 
    9.93314569703844, 10.6930904704334, 10.4763302019029, 10.6282819194525, 
    10.687132738831, 10.3998209969377, 10.4178408380566, 10.6331805354932, 
    9.30055195564525, 9.80787401101793, 9.89844269291348, 10.5207479021898, 
    9.86024499240112, 10.0318545829211, 10.6004698806152, 9.85290535308177, 
    10.2407362510709, 8.63772768159177, 9.52243374065788, 9.04652408570838, 
    8.82634645034939, 8.65287769544179, 10.1300772243523, 7.7163927936903 ;

 source_sd =
  45.6464565850607, 46.5255923443439, 51.1570028092003, 43.9613641122762, 
    48.2963987190365, 53.7611505177649, 49.1403570267233, 52.5724763487932, 
    49.2557572023189, 46.6148655024072, 51.1478387972107, 53.0637781042413, 
    63.7292570228861, 45.5412164557848, 54.7395627221586, 43.1858470587868, 
    53.1879967236506, 54.9055158728833, 46.2180793157869, 45.4582287118161, 
    40.9017370272691, 52.7964254333954, 43.774060681325, 60.2763026371489, 
    52.9834859425448, 44.7743201666019, 58.1177105922072, 58.9183153466983, 
    41.6034217716898, 41.8055263577812, 56.7807417749631, 52.9131356662825, 
    49.8340729769392, 55.6492660782917, 50.5671434540613, 51.2535394737186, 
    50.8931958538359, 49.5718166516097, 50.6890662867747, 45.0298938384701 ;

 state_variable_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 tracer_concentration_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 state_variable_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 tracer_concentration_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;
}
