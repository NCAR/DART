netcdf sgpsondewnpnC1.b1 {
dimensions:
	time = 2000 ;
	record = 275 ;
variables:
	float pres(record, time) ;
		pres:_FillValue = -9999.f ;
		pres:missing_value = -9999.f ;
		pres:resolution = 0.1f ;
		pres:valid_delta = 10.f ;
		pres:valid_max = 1100.f ;
		pres:valid_min = 0.f ;
		pres:units = "hPa" ;
		pres:long_name = "Pressure" ;
	float alt(record, time) ;
		alt:_FillValue = -9999.f ;
		alt:missing_value = -9999.f ;
		alt:units = "meters above Mean Sea Level" ;
		alt:long_name = "altitude" ;
	float tdry(record, time) ;
		tdry:_FillValue = -9999.f ;
		tdry:missing_value = -9999.f ;
		tdry:resolution = 0.1f ;
		tdry:valid_delta = 10.f ;
		tdry:valid_max = 50.f ;
		tdry:valid_min = -80.f ;
		tdry:units = "C" ;
		tdry:long_name = "Dry Bulb Temperature" ;
	float u_wind(record, time) ;
		u_wind:_FillValue = -9999.f ;
		u_wind:Calculation = "(-1.0 * sin(wind direction) * wind speed)" ;
		u_wind:missing_value = -9999.f ;
		u_wind:resolution = 0.1f ;
		u_wind:valid_max = 75.f ;
		u_wind:valid_min = -75.f ;
		u_wind:units = "m/s" ;
		u_wind:long_name = "Eastward Wind Component" ;
	float v_wind(record, time) ;
		v_wind:_FillValue = -9999.f ;
		v_wind:Calculation = "(-1.0 * cos(wind direction) * wind speed)" ;
		v_wind:missing_value = -9999.f ;
		v_wind:resolution = 0.1f ;
		v_wind:valid_max = 75.f ;
		v_wind:valid_min = -75.f ;
		v_wind:units = "m/s" ;
		v_wind:long_name = "Northward Wind Component" ;
	float qv(record, time) ;
		qv:_FillValue = -9999.f ;
		qv:long_name = "Water Vapor Mixing Ratio" ;
		qv:units = "kg/kg" ;
		qv:valid_min = 0.f ;
		qv:valid_max = 0.1f ;
		qv:missing_value = -9999.f ;
	int base_time(record) ;
		base_time:string = "15-Jul-2003,23:30:00 GMT" ;
		base_time:long_name = "Base time in Epoch" ;
		base_time:units = "seconds since 1970-1-1 0:00:00 0:00" ;
	double time_offset(record, time) ;
		time_offset:_FillValue = -9999. ;
		time_offset:missing_value = -9999.f ;
		time_offset:units = "seconds since 2003-07-15 23:30:00 0:00" ;
		time_offset:long_name = "Time offset from base_time" ;

// global attributes:
		:notes = "Only the lowest 2000 measurements are kept. Any QC failures result in rejection of entire sounding" ;
		:history = "Created by Josh Hacker with soundings from ARM" ;
		:contents = "SGP Lamont site soundings for BAMEX period" ;
		:creation_date = "Fri Dec  2 12:21:09 MST 2005" ;
}
