netcdf time3 {

dimensions:
level = 3;
lat = 4;
lon = 5;
time = UNLIMITED;

variables:

int A(level);
A:units = "meters";

float time(time);
time:units = "days";

//global attributes:

:title = "time3";

data:
A = 1, 2, 3 ;
time = 1.5 ;

}
