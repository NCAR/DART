netcdf model_restart {
dimensions:
//	time = UNLIMITED ; 
	t = 5 ;	
	lat = 5 ;
	lon = 5 ;
variables:
		
	double time(t) ;
	//time:calendar = "none" ;
	//time:units = "days" ;		
	
	double temp(t, lat, lon);
	temp:units = "celsius" ;
	
	double lat(lat);
	lat:units = "degrees north";
	
	double lon(lon);
	lon:units = "degrees east";
// global attribute
	:title = "garbage lat long for pathological model" ;
	
data:

	time = 0, 1, 2, 3, 4 ;	
	temp = 71.22, 72.314, 73.8872, 10.22, -4.222 ;
	lat = 0, 30, 60, 90, 120 ;
	lon = 0, 60, 120, 180, 240 ;
	//lon = 1, 2, 3 ;	
	//lat = 8, 9, 10 ;
	//lon = 1, 2, 3, 4, 5, 6, 7 ;

}
