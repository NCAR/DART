netcdf sgpsirsE13.b1 {
dimensions:
	time = UNLIMITED ; // (108000 currently)
variables:
	int base_time ;
		base_time:string = "1-May-2003,23:07:00 GMT" ;
		base_time:long_name = "Base time in Epoch" ;
		base_time:units = "seconds since 1970-1-1 0:00:00 0:00" ;
	double time_offset(time) ;
		time_offset:long_name = "Time offset from base_time" ;
		time_offset:units = "seconds since 2003-05-01 23:07:00 0:00" ;
	float up_long_hemisp(time) ;
		up_long_hemisp:long_name = "Upwelling Longwave Hemispheric Irradiance, Pyrgeometer" ;
		up_long_hemisp:units = "W/m^2" ;
		up_long_hemisp:resolution = 0.1f ;
		up_long_hemisp:missing_value = -9999.f ;
		up_long_hemisp:ventilation_status = "Unventilated" ;
		up_long_hemisp:height = "10 meter" ;
	float qc_up_long_hemisp(time) ;
		qc_up_long_hemisp:long_name = "Quality check results on field: Upwelling Longwave Hemispheric Irradiance, Pyrgeometer" ;
		qc_up_long_hemisp:units = "unitless" ;
		qc_up_long_hemisp:missing_value = -9999.f ;
	float down_long_hemisp_shaded(time) ;
		down_long_hemisp_shaded:long_name = "Downwelling Longwave Hemispheric Irradiance, Shaded Pyrgeometer" ;
		down_long_hemisp_shaded:units = "W/m^2" ;
		down_long_hemisp_shaded:resolution = 0.1f ;
		down_long_hemisp_shaded:missing_value = -9999.f ;
		down_long_hemisp_shaded:ventilation_status = "Ventilated" ;
	float qc_down_long_hemisp_shaded(time) ;
		qc_down_long_hemisp_shaded:long_name = "Quality check results on field: Downwelling Longwave Hemispheric Irradiance, Shaded Pyrgeometer" ;
		qc_down_long_hemisp_shaded:units = "unitless" ;
		qc_down_long_hemisp_shaded:missing_value = -9999.f ;
	float down_short_diffuse_hemisp(time) ;
		down_short_diffuse_hemisp:long_name = "Downwelling Shortwave Diffuse Hemispheric Irradiance, Pyranometer" ;
		down_short_diffuse_hemisp:units = "W/m^2" ;
		down_short_diffuse_hemisp:resolution = 0.1f ;
		down_short_diffuse_hemisp:missing_value = -9999.f ;
		down_short_diffuse_hemisp:ventilation_status = "Ventilated" ;
	float qc_down_short_diffuse_hemisp(time) ;
		qc_down_short_diffuse_hemisp:long_name = "Quality check results on field: Downwelling Shortwave Diffuse Hemispheric Irradiance, Pyranometer" ;
		qc_down_short_diffuse_hemisp:units = "unitless" ;
		qc_down_short_diffuse_hemisp:missing_value = -9999.f ;
	float up_short_hemisp(time) ;
		up_short_hemisp:long_name = "Upwelling Shortwave Hemispheric Irradiance, Pyranometer" ;
		up_short_hemisp:units = "W/m^2" ;
		up_short_hemisp:resolution = 0.1f ;
		up_short_hemisp:missing_value = -9999.f ;
		up_short_hemisp:ventilation_status = "Unventilated" ;
		up_short_hemisp:height = "10 meter" ;
	float short_direct_normal(time) ;
		short_direct_normal:long_name = "Shortwave Direct Normal Irradiance, Pyrheliometer" ;
		short_direct_normal:units = "W/m^2" ;
		short_direct_normal:resolution = 0.1f ;
		short_direct_normal:missing_value = -9999.f ;
	float qc_short_direct_normal(time) ;
		qc_short_direct_normal:long_name = "Quality check results on field: Shortwave Direct Normal Irradiance, Pyrheliometer" ;
		qc_short_direct_normal:units = "unitless" ;
		qc_short_direct_normal:missing_value = -9999.f ;
	float down_short_hemisp(time) ;
		down_short_hemisp:long_name = "Downwelling Shortwave Hemispheric Irradiance, Pyranometer" ;
		down_short_hemisp:units = "W/m^2" ;
		down_short_hemisp:resolution = 0.1f ;
		down_short_hemisp:missing_value = -9999.f ;
		down_short_hemisp:ventilation_status = "Ventilated" ;
	float qc_down_short_hemisp(time) ;
		qc_down_short_hemisp:long_name = "Quality check results on field: Downwelling Shortwave Hemispheric Irradiance, Pyranometer" ;
		qc_down_short_hemisp:units = "unitless" ;
		qc_down_short_hemisp:missing_value = -9999.f ;
	float up_long_hemisp_std(time) ;
		up_long_hemisp_std:long_name = "Upwelling Longwave Hemispheric Irradiance, Pyrgeometer, Standard Deviation" ;
		up_long_hemisp_std:units = "W/m^2" ;
		up_long_hemisp_std:resolution = 0.01f ;
		up_long_hemisp_std:missing_value = -9999.f ;
		up_long_hemisp_std:ventilation_status = "Unventilated" ;
		up_long_hemisp_std:height = "10 meter" ;
	float down_long_hemisp_shaded_std(time) ;
		down_long_hemisp_shaded_std:long_name = "Downwelling Longwave Hemispheric Irradiance, Shaded Pyrgeometer, Standard Deviation" ;
		down_long_hemisp_shaded_std:units = "W/m^2" ;
		down_long_hemisp_shaded_std:resolution = 0.01f ;
		down_long_hemisp_shaded_std:missing_value = -9999.f ;
		down_long_hemisp_shaded_std:ventilation_status = "Ventilated" ;
	float down_short_diffuse_hemisp_std(time) ;
		down_short_diffuse_hemisp_std:long_name = "Downwelling Shortwave Diffuse Hemispheric Irradiance, Pyranometer, Standard Deviation" ;
		down_short_diffuse_hemisp_std:units = "W/m^2" ;
		down_short_diffuse_hemisp_std:resolution = 0.01f ;
		down_short_diffuse_hemisp_std:missing_value = -9999.f ;
		down_short_diffuse_hemisp_std:ventilation_status = "Ventilated" ;
	float up_short_hemisp_std(time) ;
		up_short_hemisp_std:long_name = "Upwelling Shortwave Hemispheric Irradiance, Pyranometer, Standard Deviation" ;
		up_short_hemisp_std:units = "W/m^2" ;
		up_short_hemisp_std:resolution = 0.01f ;
		up_short_hemisp_std:missing_value = -9999.f ;
		up_short_hemisp_std:ventilation_status = "Unventilated" ;
		up_short_hemisp_std:height = "10 meter" ;
	float short_direct_normal_std(time) ;
		short_direct_normal_std:long_name = "Shortwave Direct Normal Irradiance, Pyrheliometer, Standard Deviation" ;
		short_direct_normal_std:units = "W/m^2" ;
		short_direct_normal_std:resolution = 0.01f ;
		short_direct_normal_std:missing_value = -9999.f ;
	float down_short_hemisp_std(time) ;
		down_short_hemisp_std:long_name = "Downwelling Shortwave Hemispheric Irradiance, Pyranometer, Standard Deviation" ;
		down_short_hemisp_std:units = "W/m^2" ;
		down_short_hemisp_std:resolution = 0.01f ;
		down_short_hemisp_std:missing_value = -9999.f ;
		down_short_hemisp_std:ventilation_status = "Ventilated" ;
	float up_long_hemisp_max(time) ;
		up_long_hemisp_max:long_name = "Upwelling Longwave Hemispheric Irradiance, Pyrgeometer, Maxima" ;
		up_long_hemisp_max:units = "W/m^2" ;
		up_long_hemisp_max:resolution = 0.1f ;
		up_long_hemisp_max:missing_value = -9999.f ;
		up_long_hemisp_max:ventilation_status = "Unventilated" ;
		up_long_hemisp_max:height = "10 meter" ;
	float down_long_hemisp_shaded_max(time) ;
		down_long_hemisp_shaded_max:long_name = "Downwelling Longwave Hemispheric Irradiance, Shaded Pyrgeometer, Maxima" ;
		down_long_hemisp_shaded_max:units = "W/m^2" ;
		down_long_hemisp_shaded_max:resolution = 0.1f ;
		down_long_hemisp_shaded_max:missing_value = -9999.f ;
		down_long_hemisp_shaded_max:ventilation_status = "Ventilated" ;
	float down_short_diffuse_hemisp_max(time) ;
		down_short_diffuse_hemisp_max:long_name = "Downwelling Shortwave Diffuse Hemispheric Irradiance, Pyranometer, Maxima" ;
		down_short_diffuse_hemisp_max:units = "W/m^2" ;
		down_short_diffuse_hemisp_max:resolution = 0.1f ;
		down_short_diffuse_hemisp_max:missing_value = -9999.f ;
		down_short_diffuse_hemisp_max:ventilation_status = "Ventilated" ;
	float up_short_hemisp_max(time) ;
		up_short_hemisp_max:long_name = "Upwelling Shortwave Hemispheric Irradiance, Pyranometer, Maxima" ;
		up_short_hemisp_max:units = "W/m^2" ;
		up_short_hemisp_max:resolution = 0.1f ;
		up_short_hemisp_max:missing_value = -9999.f ;
		up_short_hemisp_max:ventilation_status = "Unventilated" ;
		up_short_hemisp_max:height = "10 meter" ;
	float short_direct_normal_max(time) ;
		short_direct_normal_max:long_name = "Shortwave Direct Normal Irradiance, Pyrheliometer, Maxima" ;
		short_direct_normal_max:units = "W/m^2" ;
		short_direct_normal_max:resolution = 0.1f ;
		short_direct_normal_max:missing_value = -9999.f ;
	float down_short_hemisp_max(time) ;
		down_short_hemisp_max:long_name = "Downwelling Shortwave Hemispheric Irradiance, Pyranometer, Maxima" ;
		down_short_hemisp_max:units = "W/m^2" ;
		down_short_hemisp_max:resolution = 0.1f ;
		down_short_hemisp_max:missing_value = -9999.f ;
		down_short_hemisp_max:ventilation_status = "Ventilated" ;
	float up_long_hemisp_min(time) ;
		up_long_hemisp_min:long_name = "Upwelling Longwave Hemispheric Irradiance, Pyrgeometer, Minima" ;
		up_long_hemisp_min:units = "W/m^2" ;
		up_long_hemisp_min:resolution = 0.1f ;
		up_long_hemisp_min:missing_value = -9999.f ;
		up_long_hemisp_min:ventilation_status = "Unventilated" ;
		up_long_hemisp_min:height = "10 meter" ;
	float down_long_hemisp_shaded_min(time) ;
		down_long_hemisp_shaded_min:long_name = "Downwelling Longwave Hemispheric Irradiance, Shaded Pyrgeometer, Minima" ;
		down_long_hemisp_shaded_min:units = "W/m^2" ;
		down_long_hemisp_shaded_min:resolution = 0.1f ;
		down_long_hemisp_shaded_min:missing_value = -9999.f ;
		down_long_hemisp_shaded_min:ventilation_status = "Ventilated" ;
	float down_short_diffuse_hemisp_min(time) ;
		down_short_diffuse_hemisp_min:long_name = "Downwelling Shortwave Diffuse Hemispheric Irradiance, Pyranometer, Minima" ;
		down_short_diffuse_hemisp_min:units = "W/m^2" ;
		down_short_diffuse_hemisp_min:resolution = 0.1f ;
		down_short_diffuse_hemisp_min:missing_value = -9999.f ;
		down_short_diffuse_hemisp_min:ventilation_status = "Ventilated" ;
	float up_short_hemisp_min(time) ;
		up_short_hemisp_min:long_name = "Upwelling Shortwave Hemispheric Irradiance, Pyranometer, Minima" ;
		up_short_hemisp_min:units = "W/m^2" ;
		up_short_hemisp_min:resolution = 0.1f ;
		up_short_hemisp_min:missing_value = -9999.f ;
		up_short_hemisp_min:ventilation_status = "Unventilated" ;
		up_short_hemisp_min:height = "10 meter" ;
	float short_direct_normal_min(time) ;
		short_direct_normal_min:long_name = "Shortwave Direct Normal Irradiance, Pyrheliometer, Minima" ;
		short_direct_normal_min:units = "W/m^2" ;
		short_direct_normal_min:resolution = 0.1f ;
		short_direct_normal_min:missing_value = -9999.f ;
	float down_short_hemisp_min(time) ;
		down_short_hemisp_min:long_name = "Downwelling Shortwave Hemispheric Irradiance, Pyranometer, Minima" ;
		down_short_hemisp_min:units = "W/m^2" ;
		down_short_hemisp_min:resolution = 0.1f ;
		down_short_hemisp_min:missing_value = -9999.f ;
		down_short_hemisp_min:ventilation_status = "Ventilated" ;
	float vBatt(time) ;
		vBatt:long_name = "Battery Voltage" ;
		vBatt:units = "V" ;
		vBatt:resolution = 0.01f ;
		vBatt:missing_value = -9999.f ;
	float inst_up_long_dome_temp(time) ;
		inst_up_long_dome_temp:long_name = "Instantaneous Upwelling Pyrgeometer Dome Thermistor Temperature, Pyrgeometer" ;
		inst_up_long_dome_temp:units = "degrees K" ;
		inst_up_long_dome_temp:resolution = 1.e-04f ;
		inst_up_long_dome_temp:missing_value = -9999.f ;
		inst_up_long_dome_temp:ventilation_status = "Unventilated" ;
	float inst_up_long_case_temp(time) ;
		inst_up_long_case_temp:long_name = "Instantaneous Upwelling Pyrgeometer Case Thermistor Temperature, Pyrgeometer" ;
		inst_up_long_case_temp:units = "degrees K" ;
		inst_up_long_case_temp:resolution = 1.e-04f ;
		inst_up_long_case_temp:missing_value = -9999.f ;
		inst_up_long_case_temp:ventilation_status = "Unventilated" ;
	float inst_down_long_shaded_dome_temp(time) ;
		inst_down_long_shaded_dome_temp:long_name = "Instantaneous Downwelling Pyrgeometer Dome Thermistor Temperature, Shaded Pyrgeometer" ;
		inst_down_long_shaded_dome_temp:units = "degrees K" ;
		inst_down_long_shaded_dome_temp:resolution = 1.e-04f ;
		inst_down_long_shaded_dome_temp:missing_value = -9999.f ;
		inst_down_long_shaded_dome_temp:ventilation_status = "Ventilated" ;
	float inst_down_long_shaded_case_temp(time) ;
		inst_down_long_shaded_case_temp:long_name = "Instantaneous Downwelling Pyrgeometer Case Thermistor Temperature, Shaded Pyrgeometer" ;
		inst_down_long_shaded_case_temp:units = "degrees K" ;
		inst_down_long_shaded_case_temp:resolution = 1.e-04f ;
		inst_down_long_shaded_case_temp:missing_value = -9999.f ;
		inst_down_long_shaded_case_temp:ventilation_status = "Ventilated" ;
	float up_long_netir(time) ;
		up_long_netir:long_name = "Upwelling Longwave Hemispheric Net Infrared" ;
		up_long_netir:units = "W/m^2" ;
		up_long_netir:resolution = 0.01f ;
		up_long_netir:missing_value = -9999.f ;
	float down_long_netir(time) ;
		down_long_netir:long_name = "Downwelling Longwave Hemispheric Net Infrared" ;
		down_long_netir:units = "W/m^2" ;
		down_long_netir:resolution = 0.01f ;
		down_long_netir:missing_value = -9999.f ;
	float lat ;
		lat:long_name = "north latitude" ;
		lat:units = "degrees" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
	float lon ;
		lon:long_name = "east longitude" ;
		lon:units = "degrees" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
	float alt ;
		alt:long_name = "altitude" ;
		alt:units = "meters above Mean Sea Level" ;
	int base_time_spread(time) ;
		base_time_spread:_FillValue = -999 ;
		base_time_spread:units = "seconds since 1970-1-1 0:00:00 0:00" ;
		base_time_spread:long_name = "Base time in Epoch" ;
		base_time_spread:string = "1-May-2003,23:07:00 GMT" ;
	double time(time) ;
		time:units = "seconds since 1970/01/01 00:00:00.00" ;
		time:long_name = "UNIX time" ;

// global attributes:
		:ingest_software = " sirs_ingest.c,v 6.9 2003/04/14 23:15:47 gaustad process-ingest-sirs_ingest-7.5-0 $" ;
		:proc_level = "b1" ;
		:input_source = "sirs13:/data/collection/sgp/sgpsirsE13.00/1051830420.icm" ;
		:site_id = "sgp" ;
		:facility_id = "E13 : Lamont_CF1" ;
		:comment = " " ;
		:resolution_description = "The resolution field attributes refer to the number of significant\n",
    "digits relative to the decimal point that should be used in\n",
    "calculations.  Using fewer digits might result in greater uncertainty;\n",
    "using a larger number of digits should have no effect and thus is\n",
    "unnecessary.  However, analyses based on differences in values with\n",
    "a larger number of significant digits than indicated could lead to\n",
    "erroneous results or misleading scientific conclusions.\n",
    "\n",
    "resolution for lat= 0.001\n",
    "resolution for lon = 0.001\n",
    "resolution for alt = 1" ;
		:qc_method = "DQMS" ;
		:averaging_int = "60 seconds" ;
		:sample_int = "2 seconds" ;
		:serial_number = "PIR-UIR:       30682F3\n",
    "PIR-DIR:       30683F3\n",
    "Diffuse PSP:   33238F3\n",
    "PSP-US:        29608F3\n",
    "NIP:           29554E6\n",
    "PSP-DS:        30799F3\n",
    "" ;
		:calib_coeff = "PIR-UIR:     254.45 W/(m^2*mV)\n",
    "PIR-DIR:     263.85 W/(m^2*mV)\n",
    "Diffuse PSP: 109.28 W/(m^2*mV)\n",
    "PSP-US:      125.97 W/(m^2*mV)\n",
    "NIP:         123.30 W/(m^2*mV)\n",
    "PSP-DS:      123.56 W/(m^2*mV)\n",
    "" ;
		:zeb_platform = "sgpsirsE13.b1" ;
		:history = "inspired by WRF/DART" ;
}
