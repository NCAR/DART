netcdf amsua_n19_obs_2018041500.10 {
dimensions:
	Channel = 15 ;
	Location = 10 ;
	nvars = 15 ;
	nrecs = 1 ;
variables:
	int Channel(Channel) ;
		Channel:suggested_chunk_dim = 15LL ;
	int Location(Location) ;
		Location:suggested_chunk_dim = 100LL ;
	float nrecs(nrecs) ;
		nrecs:suggested_chunk_dim = 100LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nrecs = 1 ;
		:Location = 100 ;
		:satellite = "n19" ;
		:nvars = 15 ;
		:date_time = 2018041500 ;
		:sensor = "amsua" ;
		:history = "Thu Aug  7 09:42:36 2025: ncks -dLocation,0,9 amsua_n19_obs_2018041500_m.nc4 amsua_n19_obs_2018041500.10.nc4" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 Channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 nrecs = 0 ;

 nvars = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

group: GsiBc {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  data:

   brightnessTemperature =
  0.1705442, -1.235322, -1.978458, -1.769793, 0.08299936, 0.9332079, 
      0.9258245, 0.2207935, 0.6825302, 0.6809483, 0.4735224, 0.1108295, 
      -0.6032848, -1.175576, 0.2732092,
  1.283855, -0.251612, -0.7284743, -1.126574, 0.463535, 1.264464, 1.285205, 
      0.3462195, 1.154226, 1.099132, 0.9408193, 0.6478799, 0.03864326, 
      -0.4589632, 0.1675519,
  1.845042, 1.075195, 0.8709721, 0.689587, 1.186455, 1.457072, 1.442711, 
      0.07910699, 1.285423, 1.202757, 1.072864, 0.8113297, 0.3099193, 
      0.0160461, 0.06700391,
  0.8273107, 0.7740596, 1.025732, 1.606733, 1.343167, 1.474022, 1.468619, 
      -0.1428137, 1.287257, 1.230332, 1.093711, 0.8099058, 0.3529296, 
      0.1322424, -1.379802,
  -1.236446, -1.40121, -0.8141135, 0.3240715, 0.3979487, 0.7956514, 
      1.040271, 0.3817466, 0.7681929, 0.7233435, 0.5487614, 0.2454452, 
      -0.1595203, -0.452406, -0.7583573,
  -1.451746, -1.604671, -0.8616021, 0.3823381, 0.4396184, 0.8076678, 
      1.091817, -0.2279106, 0.7068119, 0.5829951, 0.4582671, 0.2042198, 
      -0.1100724, -0.5125389, -0.700838,
  -1.108427, -0.8845725, -0.4397181, 0.6902531, 0.5955248, 0.8811117, 
      1.211051, -0.7313215, 0.6802229, 0.4887359, 0.4417813, 0.1845926, 
      -0.1623592, -0.4878947, -0.6936998,
  0.004058924, 0.07525492, 0.132766, 1.067167, 0.8883256, 1.134952, 
      1.354397, -1.123105, 0.8908678, 0.6929299, 0.6599406, 0.397177, 
      0.03128761, -0.2474781, -1.084268,
  1.04817, 0.9999546, 0.09474377, -0.2935962, 0.5852197, 1.130337, 
      1.324164, -1.088398, 0.8923945, 0.6328995, 0.6399952, 0.4000587, 
      -0.0342602, -0.2347462, 0.2579373,
  1.340156, 2.020065, 0.6001499, 0.4869069, 0.9220384, 1.250754, 1.450979, 
      -1.48416, 0.9317117, 0.5893652, 0.660557, 0.4458721, 0.1319184, 
      -0.2010414, -0.2141256 ;
  } // group GsiBc

group: GsiFinalObsError {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  data:

   brightnessTemperature =
  _, _, _, _, _, _, 0.2321299, 0.2500168, 0.2500067, 0.3500332, 0.4001701, 
      0.5510925, 0.8075905, 3.136678, _,
  _, _, _, _, _, 0.3302123, 0.2315836, _, 0.2500072, 0.3500358, 0.4001839, 
      0.5511814, 0.8082085, 3.147917, _,
  _, _, _, _, _, 0.2329152, 0.2300281, 0.2500032, 0.2500077, 0.3500385, 
      0.4001975, 0.5512689, 0.8088161, 3.158886, _,
  _, _, _, _, _, _, 0.2300023, _, 0.2500079, 0.350039, 0.4001999, 
      0.5512844, 0.8089234, 3.160784, _,
  36.63401, 43.27844, 32.23582, 7.318786, 1.057506, 0.2443707, 0.2300051, 
      _, 0.2500062, 0.3500306, 0.4001572, 0.5510098, 0.8070146, 3.126185, 
      50.36055,
  11.01171, 12.94155, 9.7175, 2.289774, 0.4418843, 0.237406, 0.2300042, _, 
      0.250006, 0.3500299, 0.4001533, 0.5509849, 0.8068418, 3.123074, 22.35211,
  7.346854, 8.660736, 6.638414, 1.652725, 0.4421597, 0.2319498, 0.2300027, 
      0.2500024, 0.250006, 0.35003, 0.4001538, 0.5509878, 0.8068625, 
      3.123467, 16.91724,
  10.41171, 12.93251, 9.105816, 2.366249, 0.745788, 0.2300264, 0.2300021, 
      _, 0.2500067, 0.3500335, 0.4001718, 0.5511036, 0.8076668, 3.13803, 
      18.34681,
  _, _, _, _, _, 0.2428717, 0.23024, 0.2500033, 0.2500067, 0.3500332, 
      0.4001702, 0.5510937, 0.8075988, 3.136833, _,
  5.605732, 6.804066, 4.235401, 1.290038, 0.4440519, 0.2328792, 0.2300338, 
      0.2500029, 0.2500069, 0.3500344, 0.4001763, 0.5511329, 0.8078713, 
      3.141787, 5.215078 ;
  } // group GsiFinalObsError

group: GsiHofX {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  176.7687, 174.3334, 195.1922, 214.461, 221.9126, 220.6024, 216.2201, 
      213.0971, 209.6615, 207.6245, 207.8295, 212.1449, 220.7394, 233.5807, 
      181.5459,
  201.6861, 200.8561, 212.7437, 222.7266, 224.9058, 220.6324, 215.7015, 
      212.5381, 210.5262, 209.8768, 211.6892, 216.8506, 224.9545, 236.4631, 
      205.4069,
  235.1227, 233.8395, 239.7042, 240.4036, 233.9892, 223.6163, 217.6498, 
      214.5806, 212.6444, 212.7285, 215.405, 220.9852, 228.8233, 238.8406, 
      234.9618,
  168.3528, 172.8373, 230.9744, 246.2292, 240.0121, 228.9955, 222.7963, 
      219.4905, 217.3385, 217.0104, 218.6991, 223.8062, 232.033, 241.5156, 
      232.4545,
  160.2088, 168.0054, 223.4694, 244.0771, 241.7348, 233.027, 227.5608, 
      224.3235, 220.6028, 219.3018, 220.2881, 224.9836, 233.0938, 242.1512, 
      217.5845,
  157.092, 162.8464, 222.8916, 248.4834, 246.6255, 236.4792, 228.9898, 
      223.545, 217.8723, 218.6324, 222.2945, 228.3338, 235.8731, 243.7397, 
      215.2162,
  172.2683, 164.0731, 228.8642, 257.6087, 253.9831, 238.99, 226.9764, 
      217.6271, 211.1901, 214.9771, 220.9799, 228.1783, 236.7679, 245.555, 
      234.995,
  180.6349, 167.318, 233.0535, 259.6969, 253.1293, 236.6211, 224.4798, 
      215.4747, 210.1476, 214.5724, 221.1168, 228.8433, 238.1067, 247.3034, 
      237.6207,
  272.5648, 272.9062, 272.6275, 265.3235, 253.8874, 237.0526, 225.0431, 
      215.805, 208.6228, 213.839, 221.8705, 229.8464, 239.0799, 249.3939, 
      273.099,
  277.2926, 276.5068, 276.7426, 268.8401, 256.4739, 238.0982, 224.2647, 
      212.7991, 204.2057, 211.8224, 223.0376, 233.6157, 243.8208, 252.9215, 
      279.3009 ;
  } // group GsiHofX

group: GsiHofXBc {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  176.5981, 175.5688, 197.1707, 216.2307, 221.8295, 219.6692, 215.2943, 
      212.8763, 208.979, 206.9435, 207.3559, 212.0341, 221.3427, 234.7563, 
      181.2727,
  200.4023, 201.1078, 213.4722, 223.8531, 224.4423, 219.368, 214.4163, 
      212.1918, 209.3719, 208.7777, 210.7484, 216.2027, 224.9158, 236.9221, 
      205.2394,
  233.2776, 232.7643, 238.8332, 239.714, 232.8027, 222.1592, 216.2071, 
      214.5015, 211.359, 211.5258, 214.3321, 220.1739, 228.5134, 238.8245, 
      234.8948,
  167.5255, 172.0632, 229.9487, 244.6225, 238.6689, 227.5214, 221.3277, 
      219.6333, 216.0512, 215.78, 217.6054, 222.9963, 231.6801, 241.3834, 
      233.8343,
  161.4453, 169.4066, 224.2835, 243.7531, 241.3368, 232.2314, 226.5205, 
      223.9418, 219.8347, 218.5785, 219.7393, 224.7381, 233.2533, 242.6036, 
      218.3428,
  158.5438, 164.4511, 223.7532, 248.101, 246.1858, 235.6715, 227.8979, 
      223.7729, 217.1655, 218.0494, 221.8363, 228.1296, 235.9832, 244.2523, 
      215.9171,
  173.3767, 164.9576, 229.3039, 256.9185, 253.3876, 238.1089, 225.7654, 
      218.3584, 210.5098, 214.4884, 220.5381, 227.9937, 236.9303, 246.0429, 
      235.6887,
  180.6309, 167.2427, 232.9207, 258.6297, 252.2409, 235.4861, 223.1254, 
      216.5978, 209.2567, 213.8795, 220.4569, 228.4461, 238.0754, 247.5509, 
      238.705,
  271.5166, 271.9062, 272.5327, 265.6171, 253.3021, 235.9222, 223.7189, 
      216.8934, 207.7304, 213.2061, 221.2306, 229.4463, 239.1142, 249.6287, 
      272.841,
  275.9525, 274.4868, 276.1424, 268.3532, 255.5519, 236.8475, 222.8137, 
      214.2832, 203.274, 211.233, 222.377, 233.1699, 243.6889, 253.1225, 
      279.515 ;
  } // group GsiHofXBc

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -2208988800LL ;
  		string dateTime:units = "seconds since 1970-01-01T00:00:00Z" ;
  	float height(Location) ;
  		height:_FillValue = 9.96921e+36f ;
  		string height:units = "m" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  		string latitude:units = "degrees_north" ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  		string longitude:units = "degrees_east" ;
  	float sensorAzimuthAngle(Location) ;
  		sensorAzimuthAngle:_FillValue = 9.96921e+36f ;
  		string sensorAzimuthAngle:units = "degree" ;
  	int sensorScanPosition(Location) ;
  		sensorScanPosition:_FillValue = -2147483648 ;
  		string sensorScanPosition:units = "1" ;
  	float sensorViewAngle(Location) ;
  		sensorViewAngle:_FillValue = 9.96921e+36f ;
  	float sensorZenithAngle(Location) ;
  		sensorZenithAngle:_FillValue = 9.96921e+36f ;
  		string sensorZenithAngle:units = "degree" ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  	float solarAzimuthAngle(Location) ;
  		solarAzimuthAngle:_FillValue = 9.96921e+36f ;
  		string solarAzimuthAngle:units = "degree" ;
  	float solarZenithAngle(Location) ;
  		solarZenithAngle:_FillValue = 9.96921e+36f ;
  		string solarZenithAngle:units = "degree" ;
  data:

   dateTime = 1523756161, 1523743963, 1523743885, 1523749853, 1523755811, 
      1523755667, 1523755555, 1523755515, 1523755315, 1523755067 ;

   height = 2960.832, 3120.346, 1018.717, 0, 0, 0, 0, 0, 1689.452, 1040.189 ;

   latitude = -77.81, -73.6087, -70.294, -63.5713, -56.8731, -49.056, 
      -42.5782, -39.7299, -28.3094, -13.8741 ;

   longitude = 9.4296, 26.3631, 37.4523, 27.668, 18.8232, 25.0414, 27.1671, 
      24.8129, 29.0304, 32.5682 ;

   sensorAzimuthAngle = 296.67, 149.27, 138.63, 123.83, 109.01, 103.78, 
      102.88, 104.86, 102.21, 100.33 ;

   sensorScanPosition = 8, 25, 26, 26, 19, 17, 18, 23, 23, 24 ;

   sensorViewAngle = -25.002, 31.659, 34.992, 34.992, 11.661, 4.995, 8.328, 
      24.993, 24.993, 28.326 ;

   sensorZenithAngle = -28.75, 36.7, 40.75, 40.73, 13.3, 5.69, 9.48, 28.68, 
      28.66, 32.55 ;

   sequenceNumber = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

   solarAzimuthAngle = 144.79, 180.54, 168.42, 149.73, 129.03, 118.92, 113.2, 
      113.41, 101.72, 88.68 ;

   solarZenithAngle = 109.79, 116.04, 119.01, 123.17, 123.08, 124.64, 126.45, 
      129.32, 130.09, 129.06 ;
  } // group MetaData

group: NewMetaData {
  variables:
  	float ObsError(nvars) ;
  		ObsError:_FillValue = 9.96921e+36f ;
  	int gsi_use_flag(nvars) ;
  		gsi_use_flag:_FillValue = -2147483647 ;
  	float mean_lapse_rate(nvars) ;
  		mean_lapse_rate:_FillValue = 9.96921e+36f ;
  	float sensorCentralFrequency(nvars) ;
  		sensorCentralFrequency:_FillValue = 9.96921e+36f ;
  	float sensorCentralWavenumber(nvars) ;
  		sensorCentralWavenumber:_FillValue = 9.96921e+36f ;
  	int sensorChannelNumber(nvars) ;
  		sensorChannelNumber:_FillValue = -2147483647 ;
  	int sensorPolarizationDirection(nvars) ;
  		sensorPolarizationDirection:_FillValue = -2147483647 ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   ObsError = 2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 
      0.55, 0.8, 3, 3.5 ;

   gsi_use_flag = 1, 1, 1, 1, 1, 1, -1, -1, 1, 1, 1, 1, 1, -1, 1 ;

   mean_lapse_rate = 0.431869, 0.238203, 1.49976, 3.35676, 4.39618, 4.8658, 
      4.0128, 2.85799, -0.855057, -2.44166, -3.67322, -5.41512, -7.09678, 
      -5.56014, 0.70551 ;

   sensorCentralFrequency = 23.79974, 31.4021, 50.30027, 52.80066, 53.59613, 
      54.40013, 54.93949, 55.49868, 57.29033, 57.29033, 57.29033, 57.29033, 
      57.29033, 57.29033, 89.01 ;

   sensorCentralWavenumber = 0.793874, 1.047461, 1.677836, 1.76124, 1.787774, 
      1.814593, 1.832584, 1.851237, 1.911, 1.911, 1.911, 1.911, 1.911, 1.911, 
      2.969054 ;

   sensorChannelNumber = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

   sensorPolarizationDirection = 9, 9, 9, 9, 10, 10, 9, 10, 10, 10, 10, 10, 
      10, 10, 9 ;

   variable_names = "brightnessTemperature_1", "brightnessTemperature_2", 
      "brightnessTemperature_3", "brightnessTemperature_4", 
      "brightnessTemperature_5", "brightnessTemperature_6", 
      "brightnessTemperature_7", "brightnessTemperature_8", 
      "brightnessTemperature_9", "brightnessTemperature_10", 
      "brightnessTemperature_11", "brightnessTemperature_12", 
      "brightnessTemperature_13", "brightnessTemperature_14", 
      "brightnessTemperature_15" ;
  } // group NewMetaData

group: ObsError {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  172.21, 172.39, 193.94, 213.32, 219.62, 219.04, 215, 212.42, 208.86, 
      206.81, 207.34, 212.01, 221.1, 236.4, 181.98,
  195.79, 197.21, 210.61, 220.97, 222.47, 218.98, 214.15, 211.15, 209.3, 
      208.87, 210.71, 216.16, 224.98, 235.18, 206.9,
  228.08, 229.39, 237.24, 238.68, 232.36, 222.19, 215.54, 214.08, 211.26, 
      211.52, 214.17, 220.55, 227.79, 237.34, 232.54,
  163.32, 164.6, 222.47, 243.15, 238.19, 227.72, 221.54, 218.3, 216.16, 
      215.75, 218.2, 223.3, 230.88, 239.65, 214.49,
  169.71, 180.06, 230.16, 245, 241.65, 232.13, 226.23, 222.91, 219.8, 
      218.7, 219.74, 224.39, 232.94, 241.38, 229.54,
  158.96, 163.65, 222.94, 248.42, 246.35, 235.76, 228.49, 222.69, 217.11, 
      218.05, 221.8, 227.6, 235.82, 244.24, 213.36,
  175.54, 163.47, 227.25, 257.1, 253.83, 238, 225.91, 217.91, 210.3, 
      214.41, 220.74, 227.6, 236.86, 244.28, 229.08,
  185.41, 173.59, 236.71, 259.62, 252.54, 235.61, 223.06, 215.67, 209.43, 
      213.46, 220.36, 228.41, 237.98, 246.59, 243.91,
  271.01, 270.54, 270.57, 264.45, 252.96, 236.14, 223.31, 216.97, 207.92, 
      213.07, 220.43, 229.54, 239.3, 249.28, 274.88,
  277.92, 276.39, 276.28, 268.2, 255.73, 236.98, 223.09, 214.78, 202.9, 
      210.95, 222.65, 233.61, 243.94, 251.66, 280.69 ;
  } // group ObsValue

group: PreQC {
  variables:
  	int brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = -2147483647 ;
  data:

   brightnessTemperature =
  50, 50, 50, 50, 50, 50, 0, 0, 0, 0, 0, 0, 0, 0, 50,
  51, 51, 51, 51, 51, 0, 0, -3, 0, 0, 0, 0, 0, 0, 51,
  51, 51, 51, 51, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51,
  7, 7, 7, 7, 7, 7, 0, -3, 0, 0, 0, 0, 0, 0, 7,
  0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0,
  51, 51, 51, 51, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreQC

group: RecMetaData {
  variables:
  	int sequenceNumber(nrecs) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  data:

   sequenceNumber = 999 ;
  } // group RecMetaData
}
