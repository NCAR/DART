netcdf filter_input {
dimensions:
	member = 200 ;
	metadatalength = 32 ;
	Xlocation = 36 ;
	Ylocation = 360 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double Xlocation(Xlocation) ;
		Xlocation:short_name = "loc1d" ;
		Xlocation:long_name = "location on a unit circle" ;
		Xlocation:dimension = 1 ;
		Xlocation:valid_range = 0., 1. ;

	double Ylocation(Ylocation) ;
		Xlocation:short_name = "loc1d" ;
		Ylocation:long_name = "location on a unit circle" ;
		Ylocation:dimension = 1 ;
		Ylocation:valid_range = 0., 1. ;

	double X(time, member, Xlocation) ;
		X:long_name = "slow variables X" ;

	double Y(time, member, Ylocation) ;
		Y:long_name = "fast variables Y" ;

	double X_priorinf_mean(time, Xlocation) ;
		X_priorinf_mean:long_name = "prior inflation value" ;
     
	double X_priorinf_sd(time, Xlocation) ;
		X_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double Y_priorinf_mean(time, Ylocation) ;
		Y_priorinf_mean:long_name = "prior inflation value" ;
     
	double Y_priorinf_sd(time, Ylocation) ;
		Y_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
                time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		time:units = "days since 0000-01-01 00:00:00" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "no calendar" ;
                advance_to_time:month_lengths = 31,28,31,30,31,30,31,31,30,31,30,31 ;
		advance_to_time:units = "days since 0000-01-01 00:00:00" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id$" ;
		:model = "Lorenz_96_2scale" ;
		:model_delta_t = 0.005 ;
		:model_coupling_b = 10. ;
		:model_coupling_c = 10. ;
		:model_coupling_h = 1. ;
		:model_forcing = 15. ;
                :history = "identical to r747 (circa June 2004)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80",
  "ensemble member     81",
  "ensemble member     82",
  "ensemble member     83",
  "ensemble member     84",
  "ensemble member     85",
  "ensemble member     86",
  "ensemble member     87",
  "ensemble member     88",
  "ensemble member     89",
  "ensemble member     90",
  "ensemble member     91",
  "ensemble member     92",
  "ensemble member     93",
  "ensemble member     94",
  "ensemble member     95",
  "ensemble member     96",
  "ensemble member     97",
  "ensemble member     98",
  "ensemble member     99",
  "ensemble member    100",
  "ensemble member    101",
  "ensemble member    102",
  "ensemble member    103",
  "ensemble member    104",
  "ensemble member    105",
  "ensemble member    106",
  "ensemble member    107",
  "ensemble member    108",
  "ensemble member    109",
  "ensemble member    110",
  "ensemble member    111",
  "ensemble member    112",
  "ensemble member    113",
  "ensemble member    114",
  "ensemble member    115",
  "ensemble member    116",
  "ensemble member    117",
  "ensemble member    118",
  "ensemble member    119",
  "ensemble member    120",
  "ensemble member    121",
  "ensemble member    122",
  "ensemble member    123",
  "ensemble member    124",
  "ensemble member    125",
  "ensemble member    126",
  "ensemble member    127",
  "ensemble member    128",
  "ensemble member    129",
  "ensemble member    130",
  "ensemble member    131",
  "ensemble member    132",
  "ensemble member    133",
  "ensemble member    134",
  "ensemble member    135",
  "ensemble member    136",
  "ensemble member    137",
  "ensemble member    138",
  "ensemble member    139",
  "ensemble member    140",
  "ensemble member    141",
  "ensemble member    142",
  "ensemble member    143",
  "ensemble member    144",
  "ensemble member    145",
  "ensemble member    146",
  "ensemble member    147",
  "ensemble member    148",
  "ensemble member    149",
  "ensemble member    150",
  "ensemble member    151",
  "ensemble member    152",
  "ensemble member    153",
  "ensemble member    154",
  "ensemble member    155",
  "ensemble member    156",
  "ensemble member    157",
  "ensemble member    158",
  "ensemble member    159",
  "ensemble member    160",
  "ensemble member    161",
  "ensemble member    162",
  "ensemble member    163",
  "ensemble member    164",
  "ensemble member    165",
  "ensemble member    166",
  "ensemble member    167",
  "ensemble member    168",
  "ensemble member    169",
  "ensemble member    170",
  "ensemble member    171",
  "ensemble member    172",
  "ensemble member    173",
  "ensemble member    174",
  "ensemble member    175",
  "ensemble member    176",
  "ensemble member    177",
  "ensemble member    178",
  "ensemble member    179",
  "ensemble member    180",
  "ensemble member    181",
  "ensemble member    182",
  "ensemble member    183",
  "ensemble member    184",
  "ensemble member    185",
  "ensemble member    186",
  "ensemble member    187",
  "ensemble member    188",
  "ensemble member    189",
  "ensemble member    190",
  "ensemble member    191",
  "ensemble member    192",
  "ensemble member    193",
  "ensemble member    194",
  "ensemble member    195",
  "ensemble member    196",
  "ensemble member    197",
  "ensemble member    198",
  "ensemble member    199",
  "ensemble member    200" ;

 Xlocation = 0, 0.0277777777777778, 0.0555555555555556, 0.0833333333333333, 
    0.111111111111111, 0.138888888888889, 0.166666666666667, 
    0.194444444444444, 0.222222222222222, 0.25, 0.277777777777778, 
    0.305555555555556, 0.333333333333333, 0.361111111111111, 
    0.388888888888889, 0.416666666666667, 0.444444444444444, 
    0.472222222222222, 0.5, 0.527777777777778, 0.555555555555556, 
    0.583333333333333, 0.611111111111111, 0.638888888888889, 
    0.666666666666667, 0.694444444444444, 0.722222222222222, 0.75, 
    0.777777777777778, 0.805555555555556, 0.833333333333333, 
    0.861111111111111, 0.888888888888889, 0.916666666666667, 
    0.944444444444444, 0.972222222222222 ;

 Ylocation = 0, 0.00277777777777778, 0.00555555555555556, 
    0.00833333333333333, 0.0111111111111111, 0.0138888888888889, 
    0.0166666666666667, 0.0194444444444444, 0.0222222222222222, 0.025, 
    0.0277777777777778, 0.0305555555555556, 0.0333333333333333, 
    0.0361111111111111, 0.0388888888888889, 0.0416666666666667, 
    0.0444444444444444, 0.0472222222222222, 0.05, 0.0527777777777778, 
    0.0555555555555556, 0.0583333333333333, 0.0611111111111111, 
    0.0638888888888889, 0.0666666666666667, 0.0694444444444444, 
    0.0722222222222222, 0.075, 0.0777777777777778, 0.0805555555555556, 
    0.0833333333333333, 0.0861111111111111, 0.0888888888888889, 
    0.0916666666666667, 0.0944444444444444, 0.0972222222222222, 0.1, 
    0.102777777777778, 0.105555555555556, 0.108333333333333, 
    0.111111111111111, 0.113888888888889, 0.116666666666667, 
    0.119444444444444, 0.122222222222222, 0.125, 0.127777777777778, 
    0.130555555555556, 0.133333333333333, 0.136111111111111, 
    0.138888888888889, 0.141666666666667, 0.144444444444444, 
    0.147222222222222, 0.15, 0.152777777777778, 0.155555555555556, 
    0.158333333333333, 0.161111111111111, 0.163888888888889, 
    0.166666666666667, 0.169444444444444, 0.172222222222222, 0.175, 
    0.177777777777778, 0.180555555555556, 0.183333333333333, 
    0.186111111111111, 0.188888888888889, 0.191666666666667, 
    0.194444444444444, 0.197222222222222, 0.2, 0.202777777777778, 
    0.205555555555556, 0.208333333333333, 0.211111111111111, 
    0.213888888888889, 0.216666666666667, 0.219444444444444, 
    0.222222222222222, 0.225, 0.227777777777778, 0.230555555555556, 
    0.233333333333333, 0.236111111111111, 0.238888888888889, 
    0.241666666666667, 0.244444444444444, 0.247222222222222, 0.25, 
    0.252777777777778, 0.255555555555556, 0.258333333333333, 
    0.261111111111111, 0.263888888888889, 0.266666666666667, 
    0.269444444444444, 0.272222222222222, 0.275, 0.277777777777778, 
    0.280555555555556, 0.283333333333333, 0.286111111111111, 
    0.288888888888889, 0.291666666666667, 0.294444444444444, 
    0.297222222222222, 0.3, 0.302777777777778, 0.305555555555556, 
    0.308333333333333, 0.311111111111111, 0.313888888888889, 
    0.316666666666667, 0.319444444444444, 0.322222222222222, 0.325, 
    0.327777777777778, 0.330555555555556, 0.333333333333333, 
    0.336111111111111, 0.338888888888889, 0.341666666666667, 
    0.344444444444444, 0.347222222222222, 0.35, 0.352777777777778, 
    0.355555555555556, 0.358333333333333, 0.361111111111111, 
    0.363888888888889, 0.366666666666667, 0.369444444444444, 
    0.372222222222222, 0.375, 0.377777777777778, 0.380555555555556, 
    0.383333333333333, 0.386111111111111, 0.388888888888889, 
    0.391666666666667, 0.394444444444444, 0.397222222222222, 0.4, 
    0.402777777777778, 0.405555555555556, 0.408333333333333, 
    0.411111111111111, 0.413888888888889, 0.416666666666667, 
    0.419444444444444, 0.422222222222222, 0.425, 0.427777777777778, 
    0.430555555555556, 0.433333333333333, 0.436111111111111, 
    0.438888888888889, 0.441666666666667, 0.444444444444444, 
    0.447222222222222, 0.45, 0.452777777777778, 0.455555555555556, 
    0.458333333333333, 0.461111111111111, 0.463888888888889, 
    0.466666666666667, 0.469444444444444, 0.472222222222222, 0.475, 
    0.477777777777778, 0.480555555555556, 0.483333333333333, 
    0.486111111111111, 0.488888888888889, 0.491666666666667, 
    0.494444444444444, 0.497222222222222, 0.5, 0.502777777777778, 
    0.505555555555556, 0.508333333333333, 0.511111111111111, 
    0.513888888888889, 0.516666666666667, 0.519444444444444, 
    0.522222222222222, 0.525, 0.527777777777778, 0.530555555555556, 
    0.533333333333333, 0.536111111111111, 0.538888888888889, 
    0.541666666666667, 0.544444444444444, 0.547222222222222, 0.55, 
    0.552777777777778, 0.555555555555556, 0.558333333333333, 
    0.561111111111111, 0.563888888888889, 0.566666666666667, 
    0.569444444444444, 0.572222222222222, 0.575, 0.577777777777778, 
    0.580555555555556, 0.583333333333333, 0.586111111111111, 
    0.588888888888889, 0.591666666666667, 0.594444444444444, 
    0.597222222222222, 0.6, 0.602777777777778, 0.605555555555556, 
    0.608333333333333, 0.611111111111111, 0.613888888888889, 
    0.616666666666667, 0.619444444444444, 0.622222222222222, 0.625, 
    0.627777777777778, 0.630555555555556, 0.633333333333333, 
    0.636111111111111, 0.638888888888889, 0.641666666666667, 
    0.644444444444444, 0.647222222222222, 0.65, 0.652777777777778, 
    0.655555555555556, 0.658333333333333, 0.661111111111111, 
    0.663888888888889, 0.666666666666667, 0.669444444444444, 
    0.672222222222222, 0.675, 0.677777777777778, 0.680555555555556, 
    0.683333333333333, 0.686111111111111, 0.688888888888889, 
    0.691666666666667, 0.694444444444444, 0.697222222222222, 0.7, 
    0.702777777777778, 0.705555555555556, 0.708333333333333, 
    0.711111111111111, 0.713888888888889, 0.716666666666667, 
    0.719444444444444, 0.722222222222222, 0.725, 0.727777777777778, 
    0.730555555555556, 0.733333333333333, 0.736111111111111, 
    0.738888888888889, 0.741666666666667, 0.744444444444444, 
    0.747222222222222, 0.75, 0.752777777777778, 0.755555555555556, 
    0.758333333333333, 0.761111111111111, 0.763888888888889, 
    0.766666666666667, 0.769444444444444, 0.772222222222222, 0.775, 
    0.777777777777778, 0.780555555555556, 0.783333333333333, 
    0.786111111111111, 0.788888888888889, 0.791666666666667, 
    0.794444444444444, 0.797222222222222, 0.8, 0.802777777777778, 
    0.805555555555556, 0.808333333333333, 0.811111111111111, 
    0.813888888888889, 0.816666666666667, 0.819444444444444, 
    0.822222222222222, 0.825, 0.827777777777778, 0.830555555555556, 
    0.833333333333333, 0.836111111111111, 0.838888888888889, 
    0.841666666666667, 0.844444444444444, 0.847222222222222, 0.85, 
    0.852777777777778, 0.855555555555556, 0.858333333333333, 
    0.861111111111111, 0.863888888888889, 0.866666666666667, 
    0.869444444444444, 0.872222222222222, 0.875, 0.877777777777778, 
    0.880555555555556, 0.883333333333333, 0.886111111111111, 
    0.888888888888889, 0.891666666666667, 0.894444444444444, 
    0.897222222222222, 0.9, 0.902777777777778, 0.905555555555556, 
    0.908333333333333, 0.911111111111111, 0.913888888888889, 
    0.916666666666667, 0.919444444444444, 0.922222222222222, 0.925, 
    0.927777777777778, 0.930555555555556, 0.933333333333333, 
    0.936111111111111, 0.938888888888889, 0.941666666666667, 
    0.944444444444444, 0.947222222222222, 0.95, 0.952777777777778, 
    0.955555555555556, 0.958333333333333, 0.961111111111111, 
    0.963888888888889, 0.966666666666667, 0.969444444444444, 
    0.972222222222222, 0.975, 0.977777777777778, 0.980555555555556, 
    0.983333333333333, 0.986111111111111, 0.988888888888889, 
    0.991666666666667, 0.994444444444444, 0.997222222222222 ;


 X =
  0.323122053068933, 4.11235925990289, 10.495403938452, -1.12174943733922, 
    -1.05556850001779, 0.769627704041992, 1.8895625117467, 6.90447695677717, 
    8.68599890116947, -1.72068048915006, 3.93653221528927, 2.56087733470623, 
    -0.163502852859153, 2.62867857972446, 8.40993332089648, 1.42811357337004, 
    -3.376372206161, 0.743109048941109, 6.2870040933062, 8.84891800653066, 
    0.361024364040991, 5.14478927780334, 3.82829543195071, 0.614483196284906, 
    3.13969320018116, 6.56895575279687, -1.29194795640191, 3.14189504126654, 
    2.44685103087499, 7.94154932232449, 0.342201338521367, -3.04008775614849, 
    1.54487323459251, 7.00977637248407, 4.93037819205433, -0.871746268388839,
  8.63670835847754, -3.74913452971576, -0.685642100124471, 0.993904279720333, 
    2.28155203347724, 3.18495731856159, 6.13048014313937, 6.43680862102728, 
    -0.964475529186409, 2.42943418899137, 7.17456844496142, 
    0.276446429800959, -3.62804711545291, 0.074947570612061, 10.249439262049, 
    5.47699642685256, 0.838092443080737, 4.2369547701025, -0.274219906509572, 
    0.157641033738223, 2.53333278296865, 8.77602553233763, 
    -0.604740546812654, -1.74963308583, 0.666527989157009, 6.15227178887788, 
    5.56881003110772, -3.33697105394156, 4.56410116651521, 3.68880565844292, 
    2.77852109392236, 5.42193814547125, 3.11259922940409, -2.3278100248688, 
    1.37748020620834, 2.93484787564249,
  11.6563960425298, -2.05121057663027, -1.01533408388981, 2.67031335544902, 
    8.87340723444097, 6.1250594309492, 1.73418989886763, 3.3129808236036, 
    5.41691259027859, 0.969875369796239, -0.132010059364169, 
    4.03993043324068, 12.6015226642139, 0.667095016833629, -1.50540554255715, 
    1.68995884208618, 2.87255179496464, 4.94279096436484, -0.871967207442427, 
    -0.764773668373385, 0.779060316134024, 6.69728685792745, 
    11.2191451603935, 1.27315157170345, -1.23151834061784, 1.99404465334087, 
    9.0617514554073, 9.2248609106305, -0.363816152357486, 4.44464318500414, 
    4.66743972960976, 2.18640135842595, 5.26499181132859, 1.49505636492098, 
    0.0198111923222948, 2.50738600305631,
  -1.02714178857081, 4.59373463136646, 6.42054866158001, 0.0253863181633447, 
    3.91383538465681, 8.38167198795405, -2.33572759153147, -1.56110464365174, 
    0.176428430924508, 7.48470134797278, 1.47649701407276, -0.26161837283203, 
    2.74016273032134, 9.39504840023731, 2.07464399818244, 3.46659588068136, 
    7.29834409686209, 2.4408437574241, -4.12044692163553, -0.225711438713845, 
    2.69575708165322, 9.04650272309986, 2.7326425448002, -2.25775118814345, 
    -1.2990123263732, 0.150611134016191, 2.461631552588, 4.29833261559302, 
    6.8536853348101, -1.99711799412616, -2.07269151990527, 
    -0.410455844162249, 9.95744667379301, -1.5803810797941, 
    -0.10775247627181, -0.973085783126263,
  1.27586636316947, 2.5315591180758, 4.44503787978176, 5.04093946023139, 
    0.964092142369453, -2.47142793445914, 1.5980493816187, 7.27682158861053, 
    9.91608628782452, 1.46676968547661, -1.16709815598815, 2.55613863731139, 
    8.70497683482648, 5.49966538895321, 0.622253106323619, 4.82119128300163, 
    2.23186111135668, -1.05967172101883, 1.91591265275321, 7.01200783430546, 
    2.13036503703981, -3.45334803427381, 1.94529739845056, 6.77525777242481, 
    3.95001543087835, -3.36979214328696, 2.69932963065762, 3.71092469700676, 
    5.78829479118628, 4.23026146705175, -1.7210953318297, 4.14071040561375, 
    6.30698433471232, 5.4423223267915, 3.79302134621202, -3.52305422451557,
  -0.380789243856788, 0.733036940264083, 2.95013699922518, 8.79387214322292, 
    -3.35057891063328, -3.15110323631558, -1.50946989587164, 
    6.99312038601452, 0.427675532368032, -2.31174648756589, 1.57357161627712, 
    5.95361254027035, 8.23485620517622, 1.49184422192118, -3.99803362638296, 
    1.18325544649512, 0.684967297844757, 1.78357317965209, 3.49609295126671, 
    8.29535049154808, 8.30179422533367, -3.19886244564514, 2.19564270334191, 
    6.00900086687881, 5.55396291455208, 6.02610726799593, 5.33918878174608, 
    -4.65354780199958, 0.528537104400728, 3.62733738727574, 8.91928213362464, 
    1.27766067836919, 3.80139412484568, 7.70652452389342, 2.12169359610505, 
    -1.77514002482177,
  3.59019796045997, 1.87812618914157, 5.107120101615, 8.30009064585059, 
    1.85950370007138, 0.508904996109866, 0.101563400219494, 
    -0.458140327632194, 1.65468114379677, 7.40671131588429, 3.09399761735785, 
    -3.667525992281, -0.270757380923831, 0.892359055381582, 2.69376484642959, 
    6.11255520034459, 4.67811049520342, -3.75204451081345, 1.65125175189989, 
    2.74315952640067, 2.54285675334064, 4.57752850415818, 8.33228851560077, 
    -1.59129799730938, -2.87458566295544, 0.00405310598975817, 
    7.53823966428021, 2.01967164311791, -2.46318985729916, 6.00832972059579, 
    4.60381991698812, 0.898892980173189, 5.46603830542342, 10.5822445502718, 
    -0.90709708864658, 3.15758678510373,
  4.55655261045657, 8.31218805246818, 5.08922846950804, 3.7032477519865, 
    -0.83282780939355, 1.87272912050023, 6.33950594305644, 4.99826991641584, 
    -3.48540881685002, 2.32327999862117, 2.8742702817551, 5.83828432806283, 
    4.48340544286193, -3.87928703999689, 2.86127917437242, 1.90484757670062, 
    2.23482438285232, 4.7066660742142, 5.73881094776736, -2.56130685468527, 
    -1.39732912820109, 0.886185590460258, 8.05537517842535, 5.0684432908533, 
    -1.7679968842981, -0.32668114207728, 0.370289981807412, 2.95682733150687, 
    8.29064879536328, -1.37460624102255, -0.858666130650466, 
    0.560092084359741, 2.56338644550987, 6.74129268691379, 3.56652745844778, 
    -1.38435903784728,
  3.03100826592502, 5.01668381694902, 5.81575900521723, -2.62098703809075, 
    0.940020192970306, 3.63319851682718, 8.60601129754569, 
    -0.770911907222531, 3.29424358741393, 2.45597463778315, 3.51048714383034, 
    6.53543037443353, -3.78670307605664, -1.70763878142069, 
    -1.41936539624014, 5.13161099139387, 8.96890154484881, -1.43156480731205, 
    -0.301833704523819, -0.950763765992303, 0.845161897459062, 
    2.66030837905816, 5.75719411997133, 5.11166307666213, -2.53943212663568, 
    0.696224800180287, 3.04043356514238, 8.31219727050601, -1.9517650882823, 
    2.89434156540051, 2.51049231327806, 5.18741771121538, 7.69708955806104, 
    -2.19385261051543, 3.52560537891954, 3.79027202843235,
  -1.16563273901807, -0.34699291937274, 8.80401474979293, 0.691166571345053, 
    -2.65291284415414, 4.47121444129705, 6.84242846381339, -2.35659252518696, 
    2.31911763966548, 8.4676580763238, -4.04655524382492, -2.96356900309089, 
    -1.49944352338795, 7.43272394055584, 7.40499478989827, 0.198527566440734, 
    1.75535754225472, 4.56665715197527, 6.37873289134237, -1.78549589277698, 
    -1.5450841455467, 2.00962296116361, 9.87921650086772, 4.70358876525971, 
    2.47669816980005, 2.68598346578885, -1.83477346195018, 0.945971075981722, 
    2.04747886313724, 4.66851763262538, 6.28570260479404, -1.68839748966612, 
    -1.38721624498427, 0.912904176918421, 9.49511628447865, -1.72182663007112,
  -1.0177248551582, 0.614662217932558, 5.28522929561208, 3.59854807107019, 
    -3.84349950633411, 2.46086534922287, 3.17003999416116, 6.84290321216625, 
    9.15099212167934, 0.915625874141745, 2.79842396774192, 2.4548229727208, 
    -1.4337567844023, 2.87755410096288, 4.41504004589541, 5.10780200593065, 
    5.34731011676944, -0.647287399822243, 3.27972173914133, 6.33204694939101, 
    3.15332956959356, -3.03588786579556, -0.689937734289168, 
    1.09860981682699, 6.87011222547555, 3.77266797723587, -2.36742769793655, 
    -0.511757193886621, 2.3655276545511, 8.07567741275984, 
    -0.728605994501999, -1.9042643503923, 1.63994607908307, 6.03972810248243, 
    5.62322923654374, -3.06800930552353,
  -3.16179455172978, 0.232763838101207, 1.20016017619631, 8.21972546379374, 
    3.21316013671926, -5.91635607389969, 1.07085640206026, 
    0.0696855798466709, 7.07220276707807, 1.92243186087521, 
    -0.246877665835206, 2.37598487058803, 9.555165009477, -0.372285575506373, 
    3.86480637995857, 1.78478818686483, 1.86559754364566, 6.99295317652549, 
    6.41285893289839, -2.75207265302132, 2.55949078758473, 1.76112178048951, 
    1.55343024641683, 3.35332057009633, 6.08281988632263, 0.265969095067391, 
    -2.79803237906373, 1.28959223144627, 3.31230420074055, 6.78249383897736, 
    0.226804005312647, -3.03088931728292, 1.28491387192532, 3.14559875917784, 
    5.61468352581143, 3.47368817442179,
  4.28504865203381, 8.01528605060255, 0.798838588797347, 1.80046057472189, 
    5.5279366366749, 4.5553706148719, -2.87943058698482, 3.29810838941007, 
    5.24750083553265, 6.4049567693135, -4.28164358111204, -0.117265085945767, 
    -1.36276209891543, 7.98593799240956, 7.34093689721586, 2.38460631688237, 
    4.18485378403743, -2.94363533162073, 0.628886103242686, 0.96523170418673, 
    2.7840566418676, 5.2721715581102, 5.22725671041108, -0.852447652028598, 
    -2.03569040847709, 2.23051546740201, 7.04341735494565, 5.25249710923659, 
    -0.340968692263347, 0.587218896970955, 5.95602053701695, 
    9.32729754140691, 1.07066024588818, 1.96671869472852, -0.732732855138443, 
    2.12168931874095,
  5.58481070903527, 4.37321927580485, 2.36180631360739, -0.682033069157917, 
    -1.55845092471456, 1.04603316836454, 7.59778640196042, 3.69064507755884, 
    -3.25530981650432, -2.31436183626479, 1.38515769730442, 3.97809736161642, 
    6.34889687756492, -0.327215325731477, -2.15316057676941, 
    1.47703097522474, 10.8834613175045, 3.48543402117659, -1.04971611339381, 
    0.234127241242661, -0.474597421013999, 2.29060274614381, 
    10.0347504957409, 2.91547971517003, -0.337490563094515, 1.62269274538874, 
    1.08571208007891, 4.07389466736695, 7.66983522518106, -2.59153762995878, 
    -1.24366749035249, 0.225064627916423, 4.66114849844904, 11.6356343701163, 
    0.867282941090589, 1.57069496288443,
  -3.03557599583543, 1.04233819194959, 2.15226481609975, 3.3057990115052, 
    5.43705208904772, 4.86486969300509, -3.22008194817254, 1.15287307769732, 
    1.05016909497958, 2.836574213562, 6.62266108801036, -1.73298837431823, 
    -2.11507183475671, 1.70484695151722, 3.21857227298637, 7.33296882970679, 
    6.86223936953341, 0.436573074327732, 6.02663612223056, 3.38229695417427, 
    -0.195957997009011, 2.97989545419297, 7.31515673562356, 
    -0.230754449543966, 3.08472035951278, 4.99258010352021, 4.95381384915308, 
    -1.1447462388683, -2.8996303942587, 2.49799656422549, 7.40250609918777, 
    6.58922777768408, -0.506435893001215, 0.45025086341003, 4.30983473972981, 
    7.48742806279585,
  8.837695412513, 0.26763494840339, 3.48068374880243, 5.03310096844391, 
    5.74767776570101, 5.1035681204268, -2.53879041018707, -2.19120146409119, 
    0.916317475731251, 7.02330228437486, 5.48123404991873, 3.1091312506256, 
    2.25318010631837, -2.73588178035911, -0.524791219977382, 
    1.15385907401667, 7.30374414019316, 7.81251931444277, -1.61166825387677, 
    -1.03358204014533, 3.94670091850381, 6.86130466595466, 4.29364668080533, 
    5.08614225953435, 2.51748479246194, -0.820772800741803, 3.57339971276033, 
    8.31984582225449, -3.2543349237278, -0.402407311681398, 
    0.449475663452972, 1.44309250769211, 8.19527593971874, 
    -0.00511173509219898, -4.32844878426993, 0.64331161089736,
  0.23247442204582, 7.96473120658077, 2.33173372274518, -0.509528454625491, 
    3.46575728085867, 6.33531882336502, -3.05624940658794, 2.6488350599772, 
    3.76216173353014, 9.71780350128565, 1.90130360048832, -3.82312332603315, 
    2.12480498534171, 7.537887139209, 10.2279274875762, -2.15462940077763, 
    -4.12743488032275, 3.28303395783279, 2.93535736208304, 1.32992885006159, 
    5.08999321917718, 9.28233067757629, 2.58715149167382, 4.14089973987527, 
    5.04500290572259, -0.261589354589042, 3.49306551824573, 5.65937251603872, 
    -2.87776364427887, -0.748378145020112, 0.564073047757656, 
    2.55764781508966, 6.33888268040809, 3.63663463903565, -5.02186978826651, 
    0.911775679641784,
  4.10752801529527, 5.54524434539528, -2.98033435654244, 0.628004236436859, 
    1.38374237791025, 4.24805469178051, 4.85159796938708, -5.30238719300732, 
    1.60947910416616, -0.26940529455601, 2.57492568104719, 11.4197681132535, 
    -0.687414935570549, -0.788182999105865, 3.7036959222451, 
    7.21953080381129, 5.91784739085525, 0.305529662612122, -3.28861649883763, 
    3.41093672393041, 3.97530659246911, 1.63577827525022, 3.10745693457167, 
    7.1545402831987, -1.35159091715058, 4.19990200946202, 0.478486782445637, 
    1.94438033428688, 10.8726304739025, 6.63087107922717, 2.39323007881488, 
    4.57800263467132, -0.165060699321507, 2.78363799498923, 2.32043735222094, 
    1.93286914910427,
  8.88589097230201, 1.02367803429387, -4.66836685359793, 2.89660199643602, 
    2.64437157222636, 2.75845325636824, 7.25606730433973, 5.27936756541806, 
    -2.61438271075916, 0.386345866759648, -1.29109797586642, 
    0.843666234683775, 4.39922881383243, 8.88440058017963, 4.07449107346665, 
    -3.16088675745474, 2.55210887632793, 7.34851635027226, 5.84995581433, 
    -0.525806111480926, -2.00128973439909, -2.23843028565668, 
    -0.64159401494836, 4.62226400417708, 9.36833519212991, 2.05549662491576, 
    1.07498763751567, 2.84027627343332, -0.712876820013214, 
    0.305389970900955, 1.4673376959835, 5.79419629126913, 4.32939008830614, 
    -4.63107174341427, 1.48492465638702, 0.118715444302638,
  6.83638765182475, 8.81206060770563, 3.95385562303367, 0.440808060113397, 
    -2.21143022817581, 1.87281187137758, 1.91569162803956, 0.700624355751222, 
    1.13843353629152, 7.64268539473184, -1.0947059789289, -1.73502184786176, 
    -4.10618750193593, 9.05282331731505, 5.2569924397808, 0.609111393414459, 
    2.66857441108353, 8.79314829139701, 6.83225197930258, 2.24519817539261, 
    5.89632206859919, 3.96476440918654, -0.499657133772896, 
    0.896146440319175, 0.289877591044227, 1.91070976090902, 5.08250392739952, 
    7.49684152975657, 1.5048613197502, 0.15322603945302, 5.24595176984512, 
    10.9428749589669, -2.23106576207587, -1.59236017260016, -1.2587798951797, 
    0.698489820289734,
  -1.70402400077425, 3.04544914439609, 8.7513363927646, 3.19509875829814, 
    -1.8221603525465, -1.72645605380351, 1.86352177327253, 3.19792133690002, 
    4.41726801748568, 6.97073974635715, 0.633251682516071, -3.94477053535092, 
    0.923132047825226, 3.71463840658643, 6.85682796774068, 3.73857218597281, 
    -1.34140567259732, -1.48552212307251, 0.486339236004362, 2.0142391866138, 
    7.6204420359923, -1.04145030160769, -3.98207003378803, 1.69205738744671, 
    2.07970998448193, 8.45171505935152, 5.7690188084892, 1.38141011443817, 
    7.21702413298736, 5.07128804610836, -0.979608970491493, 5.22694374233683, 
    7.39197648750876, 1.88477450004816, 4.22992733075919, 2.44109861486746,
  0.0322310973573843, 0.589357992879836, 4.28465075832616, 6.54885864448609, 
    1.11827700679414, 3.14500928911434, 5.84453076252651, 0.500381857947761, 
    -2.36965493784557, 1.93011317726355, 5.77179573848821, 5.54249599030343, 
    -2.86725039391766, -1.38715348083749, 0.464990458652413, 4.4086995183734, 
    6.95417136344985, -2.81174152138093, 0.303267472564354, 
    0.606397433021395, 2.58850174436305, 6.96156945894087, -3.12418558948976, 
    -1.81102938227346, -0.40371390296653, 5.26217952306348, 9.69095281676302, 
    2.27232374146919, 3.64624035936104, 5.57919133149293, -1.68065851763643, 
    0.00105090590149937, 0.44540715217818, 3.31205965094949, 
    10.4341328401468, -3.36987495321511,
  1.40011225065598, 6.92806203980646, 6.61402010048013, -2.91502488994595, 
    -1.53370243392563, 1.78787700277625, 9.21805938320925, -1.93960751888874, 
    0.968989777549559, 1.66262429260049, 5.72706302975072, 4.26045334869613, 
    -4.00418678093364, 3.06653967584338, 4.84696309060713, 5.62406257425258, 
    -2.53449478463279, -0.5900809223649, 1.18544544739318, 4.06582973613876, 
    8.25782437547616, 1.43757821117727, -2.28884314462595, 3.88934345662456, 
    6.38177827667793, -1.20680968217998, 2.75029535660701, 6.0599754576593, 
    4.59672094627408, -2.90878390374015, -0.325875394430186, 
    1.19034512380313, 3.8720814261086, 6.06064349713043, -0.258207724960943, 
    -2.37800708886628,
  -0.44028964545288, -0.861926667490681, 4.13684078694189, 9.96075764814052, 
    -0.983449651547337, 1.15248290380133, -0.60978528756129, 
    1.42928202299438, 4.469754782905, 8.46284222803598, 0.61376663545643, 
    -5.59789833363223, 0.566728766348374, 6.7003518149853, 5.17154454912998, 
    5.13472772087626, 8.93325161864268, 0.385059281854461, -4.74539566974513, 
    1.59796158046433, 6.26859950352971, 1.51444082368749, 2.11963169288719, 
    3.85943384300413, 5.09479336113661, 5.99670480629373, 3.30000329167689, 
    -1.80239903380529, 0.734549087176903, 4.68159256304784, 8.68866511471497, 
    -1.85606985938138, 3.49055596641112, 3.38585342949713, 4.51449916225686, 
    7.53616998941712,
  6.56095071433369, 0.424050651995128, 4.71922591696298, 4.11403111200831, 
    -3.17895891241244, 2.8302726246323, 4.42486548908004, 5.50707167704083, 
    3.84352536970783, -2.4352147886845, 3.28222379029213, 5.67206965881073, 
    5.85262878047441, 2.46878091760565, -3.08770250827574, 1.45254342938632, 
    4.81783017373109, 8.01384533252082, -0.0050579071509933, 
    3.90658365813587, 4.45372450193588, 4.21691574779392, 4.46779895002205, 
    -1.70976929107254, -1.44805792956832, 1.01488315906889, 7.55996915253064, 
    4.52758597527808, -2.74244956330549, 0.020314970210026, 2.5348800688955, 
    8.88079982347592, -5.0264501529638, 1.37933709301126, -2.19169346138696, 
    4.30794897214674,
  4.27611120233472, 5.40501829945088, 2.80136561029305, -0.479437518443499, 
    2.91958634039849, 8.29525442931876, -0.413969650995371, 3.98595088955833, 
    3.84197487049094, 4.48776114624775, 6.21043407119966, -2.36750767488169, 
    1.23306323403231, 1.77217605789083, 6.47104021071086, 4.64747279628157, 
    -1.81510550336893, 5.57098176267956, 6.11540401420813, 3.69304816308251, 
    6.09321016711379, 1.79489330861528, -3.2873914916341, -0.303457300350851, 
    0.317248938065751, 3.72245694614039, 8.45289963680961, 
    -0.472729957012267, -2.18884739278638, 0.560615082442396, 
    1.42034540706548, 3.17884988629904, 5.77944476534797, 0.0644142050184806, 
    -3.90923344819971, 3.2221475879759,
  -0.740594078083789, 3.22065850213393, 10.5044089867963, -0.474287896720751, 
    -2.11864466672458, -0.149408261983563, 0.894968308285698, 
    5.99697972251697, 2.2536924504581, -1.73650840263104, 2.23972382788453, 
    8.34049758894491, -2.7019634870792, 0.514823413165149, 
    0.00490535201976616, 1.71971353339521, 7.92021803489685, 3.6353707231681, 
    -2.28994888398007, 0.865946661571, -0.32757045802058, 1.1911855683975, 
    6.6629089261916, 3.31280922722764, -3.4276854782437, 1.24841124248279, 
    2.3745432471925, 8.647737631436, -3.20969268135111, -2.43184147620861, 
    -2.14022583072302, 7.05307954546234, 5.95544898756303, 1.71388663303543, 
    5.66933804284517, 1.76893290176878,
  6.17448979868222, -1.49164455065633, -1.57305318308991, 1.60218460212821, 
    8.43528143205147, 6.81598516294651, -1.04875283289172, 
    -0.772085645255334, 3.7330387398966, 10.2793520650836, 1.23926819931681, 
    -0.089166292506615, 0.711086028941653, 0.0946209180735975, 
    2.91590467757505, 9.46747210280333, 0.25017545431478, -2.4066428697743, 
    -0.559775903412541, 2.72567924098125, 7.43904031604186, 5.37850600743214, 
    3.62751963197184, 2.26058710450547, -0.362139330430902, 3.06506261573468, 
    6.90378653613019, 0.642314847918678, -2.68840690928263, 
    0.897100795112878, 2.40333553847948, 6.90045223496393, 
    -0.744842933309958, -2.09426516517569, 0.904626341468107, 3.60471974791669,
  -2.16943287688458, 2.591969727168, 6.78557631301806, 8.70574245144231, 
    -3.28463265744259, 2.36332232531981, 3.33197522431844, 2.18702833691144, 
    3.66765697935932, 6.18508065499133, 3.18846557888495, -1.89347098406381, 
    -1.13337958639037, 1.36723878203273, 4.78514733184716, 6.06566369235365, 
    0.309482018478414, -2.7747483863587, 0.645146711447335, 1.89289201688796, 
    6.31021065060668, 3.5831791378882, -4.09302929676952, 1.09084577155937, 
    2.24197843275635, 5.69564741868135, 5.9784854967832, -1.98668566037263, 
    -1.09349825831267, 2.1707604551777, 9.99196100544169, -0.869347264949214, 
    -0.285396408013134, 0.92987960424033, 4.09400465435805, 7.13844738088591,
  2.00216957819037, -0.881749099659254, -1.29304230078714, 1.49176748290685, 
    5.57314061916529, 5.26748324023371, -3.24285607810871, 
    -0.317997266415712, 0.369579812991285, 6.08046289270773, 
    3.94544081090955, -3.56166598910432, 5.13493617861345, 2.69122551502827, 
    0.590664255608332, 3.47561169897863, 8.63668885899758, 0.325825346940233, 
    -1.82108687049651, 0.288921563912212, -0.178513572183911, 
    -0.717446452641784, 4.89445974468627, 5.71015008494647, 
    -4.18956213090281, 4.97667931402679, 6.0931788168351, 3.21212793018922, 
    4.95191414535431, 5.75494499532652, 2.77587081280673, -1.33422781281494, 
    -1.79061714479837, 1.42176343159674, 6.22887344316456, 6.05278066204067,
  0.663009860994316, -1.7754161022209, 1.06358999421086, 6.54805275871338, 
    6.23812873461996, 0.0183997339089355, 0.379187071355154, 
    0.641342967003214, 3.28870656178518, 2.34499407557569, 2.97303920025433, 
    2.37641644471094, -3.17948842396722, 1.63092815703388, 4.92060476416325, 
    9.72532798282689, 5.74547807534399, 4.1316544919232, 5.51515582738565, 
    -0.70889417055421, 2.67292177872009, 5.6563799501853, -1.58520439977489, 
    0.126597962462915, 2.1360615105861, 5.0428903991237, 5.69028130503868, 
    3.09961159028507, -1.43252149726755, -1.21183636371512, 2.54666115848239, 
    7.68823607460391, 9.11498942456255, 0.875123861822564, 
    -0.218184187127909, 6.83508865219304,
  1.62782358548285, 6.736312434016, 4.47904605599215, -2.47678113377192, 
    -0.460876788274185, 1.25871374443652, 8.16483851265189, 5.86856716248456, 
    -0.548064374357092, 4.80991795269159, 7.7089457958186, -1.79253235122471, 
    0.317482847873789, -0.174726345233882, -0.0326447318246506, 
    0.630645176161749, 5.58365582081142, 7.39927350840747, -2.82591617611485, 
    1.45767649736929, 5.91441838091604, 6.80418998306646, -2.97132304437209, 
    4.72040562270274, 3.45639638834108, 1.47712405954455, 3.93942203109058, 
    7.12386881276482, -2.64168293558186, -0.82324643896273, 
    0.311884323375347, 2.58373020937443, 6.0285206588552, 4.47046942225219, 
    -1.84797136650104, -1.3325020713252,
  8.00831831642528, -2.66104936256719, 3.333793696443, 5.13586516403591, 
    3.93052872872842, 4.54596222378085, 2.03690116042078, -4.29455054439392, 
    2.14760615557801, 3.02459167475264, 5.15165270880918, 5.17710913002746, 
    -2.1048326082623, 3.90954921699722, 5.33837046557992, 5.47649214252439, 
    3.66256304494216, -2.07552830912407, 4.41766947977813, 6.28871562903653, 
    4.5116378945379, 5.43217818237822, 0.722821916088972, 
    -0.00266127706366248, 4.69604665738803, 8.85505945927014, 
    0.294462735685475, 0.630729349735467, 0.00905577724439199, 
    2.62867210834212, 7.04589096833961, 3.21799498916775, -3.2970560020696, 
    -0.30604264271227, 0.813983215271285, 5.75664153218005,
  3.62680702458811, 3.05313641416114, 4.36880476181679, 8.05528101318535, 
    3.27604090758379, 3.9578740975158, 3.96746333084568, -3.79295894711139, 
    2.72118716208376, 2.94040747195173, 10.0551638365515, 1.25045725147695, 
    -1.26394328375807, 5.13909867987302, 3.84418993736347, 
    -0.0455763137252578, 2.88882063591443, 6.75731926264214, 
    -0.727693521359745, -1.90083856682299, 1.64106681593788, 
    6.38038333850267, 4.59853254255197, -1.66655083264834, -1.3319036230275, 
    1.31615543586586, 7.63573303780212, 2.73431029894169, -4.1355259959573, 
    0.802079519805061, 1.49504425981569, 1.80381795291193, 2.7862327268362, 
    5.81020672757576, 1.87775451542357, -5.93475319612889,
  2.88372512495633, 7.09072455691407, -1.85068608768144, 3.03941538620751, 
    2.67141044550617, 2.78542561701346, 6.66795363653737, 7.07390608009297, 
    -1.06771907840255, 2.60425391908991, 2.16163945567081, 0.419522527888717, 
    2.55329277483094, 7.9350265147384, -1.68621231274287, -3.84712170093331, 
    0.655539933103617, 2.81734579836178, 7.04893560380766, 1.22656867681533, 
    2.07506811372361, 3.77622076829903, 9.13023949416985, -0.728550017767248, 
    -0.50284728153882, 2.00220746141071, 10.000349382745, 0.536811583799667, 
    -1.44523478841239, 3.42423654150757, 2.67494836717753, 3.5920782485088, 
    6.59818317888975, 0.277687127348915, -2.46976465149721, 0.841832007788932,
  0.232444172617209, 9.11032048041963, 8.18134671832068, -0.279938736055289, 
    -1.73940781378166, 1.51453078355056, 1.84859859721802, 1.48968696761889, 
    4.48090486036045, 9.37210538071841, -1.89955600850414, 
    -0.434088451226301, 0.97237556729761, 0.33394994059417, 
    -0.369178760236971, 7.08366114476472, 4.9302503371521, 
    -0.451057390841733, 4.70281656795896, 10.5786660553651, 1.97286127071206, 
    4.64830138468725, 8.38474996822098, 0.244935999931771, 0.737904516159454, 
    1.35762114572545, 0.404021960480112, 2.59787215584229, 6.80711114568591, 
    -0.477681660010814, -2.8526906844592, 2.0852911468731, 3.22914588506269, 
    9.19090627266093, -2.79599578414952, -3.71556980589451,
  6.04764522256497, -2.55966102152109, -0.0142317077279479, 
    0.916809456861439, 6.0459645032503, 10.1620782585135, 3.12119872789046, 
    3.5799523463054, 3.00501818784043, -1.91106150382263, 3.92644133671657, 
    3.74134509099508, 3.20297292270299, 7.02025476280962, 3.50347829049196, 
    -3.36642336143844, 4.01763294201454, 7.05600978421071, 2.73282183785548, 
    4.57303768403174, 5.38082421469558, -3.11713552034567, 0.727231572878793, 
    1.04646388012107, 8.4216540995921, -1.27004660290936, -0.881719493971835, 
    -0.427329032052012, 10.5263543333757, 4.24637026192609, -0.9387440727747, 
    3.74076812240208, 0.461440656014957, 1.63563115251333, 2.45815825401244, 
    5.12112701354201,
  2.80863889705779, 8.4388236613799, 0.381103730292308, -2.2377329090263, 
    -0.0726728762370477, 1.26597790405041, 2.54002027247648, 7.6539956068164, 
    -0.799784597330549, -2.3088941987561, 2.62635787112759, 6.36301359468518, 
    4.23636834741063, 3.71228065055505, 0.390586067010092, -2.12401732103218, 
    1.45391982442503, 3.70924770955971, 7.14679294933874, 2.42801128806361, 
    -3.07727468446329, 1.38070201482132, 6.02036298819823, 2.27039587017949, 
    -4.72512908617665, 2.61527114780816, 4.08448001654487, 5.80991065715294, 
    6.20789401833172, -4.99193429024318, 2.40961979665617, 4.14687523367226, 
    8.00355482820712, -1.57601753071156, -0.511855971640765, 0.184735863060709,
  4.36834643088447, 5.18833760942122, -3.33539344237365, 2.08084679784347, 
    2.35560624073173, 8.27491241508533, 2.97561037765022, -4.51012167015735, 
    2.53832404730225, 7.22493586466674, -1.08681305440164, 0.219231553293576, 
    2.10978605737134, 7.8761722463044, 1.89186458622323, -3.59005470712212, 
    2.20032199626428, 8.27846306938466, 3.68469765775752, -3.33405928224638, 
    0.319244173035136, 3.72555612463769, 6.70177173505554, -1.81528050049844, 
    3.61896578190781, 6.25131558297302, 5.52040106234434, 0.985164602950922, 
    -1.29194645418973, 3.14791911362845, 8.8982327391401, 4.41836186205087, 
    -1.15631209555525, -0.892100761934346, 0.435106482701897, 1.60312696812118,
  -0.94522967224791, 4.05877073723767, 6.51750614077211, 5.80815527782957, 
    2.49317991085035, -1.12327528138394, 3.82866659294086, 9.33600856711271, 
    0.43767292089043, -2.94588901288553, -0.666347913538275, 
    3.91087381506225, 8.31124423637597, 3.06922402125145, 3.66747863431599, 
    1.89671182745222, -2.6173943988024, 1.84181340448191, 5.00445988692074, 
    6.70711746172364, 2.31977633054194, -2.02452671247957, 
    -0.562538830606109, 1.03028288754328, 3.22242849306806, 6.27176720714497, 
    -1.65520736043545, -3.26440965370861, 0.862546691767485, 
    5.22756220070046, 6.48200302340128, 0.0253886612238507, 
    -2.15964733359267, 1.32119498174615, 5.43948243632683, 6.68395497102473,
  -3.27409606335833, 3.72627166494257, 4.8740279694715, -1.66465203563221, 
    2.97319889931187, 3.78473112113607, 7.07344793061554, 9.07578914454794, 
    1.81001278367423, 4.32076394105135, 4.78761865089717, -1.30444625818336, 
    2.70762770641693, 1.76367988532528, 1.94723409359659, 4.6737016368511, 
    8.15372566958979, -4.28774712080387, -1.65840995223414, 
    -2.28921253527592, 9.28049948423053, 2.55900057946062, 
    -0.104955301536609, 6.45198937797055, 4.79419034305486, 
    -0.208071592010989, 4.24743826560398, 10.0669680964273, 1.61789250192873, 
    2.61732763966991, 5.22403183911048, -0.355813711682445, 1.05529908432082, 
    3.11480784042025, 8.94268047660495, 5.63094651727515,
  -1.18042532297014, -1.43243511696147, 1.22258185890922, 4.15922225667182, 
    7.16891544895632, 0.14810792557269, 3.11324672331054, 6.69218649414929, 
    6.77305547672086, -1.00354951831857, -2.19379183049217, 1.31966707469594, 
    8.20238851353893, 0.965309113645715, -0.301529757317688, 
    3.44681437210546, 8.65742878869533, -1.48984786258007, 1.99804635969697, 
    7.41895034026801, 7.36481791363751, -1.50991560312181, 3.83535685088006, 
    3.10768785731608, 1.05643902421968, 3.72776264215056, 6.15770938456259, 
    -2.63652414509751, 0.638485850183419, 2.12916869340959, 6.13871876664469, 
    5.92691205585797, -1.60334847298655, -2.03132855088113, 2.52054103230912, 
    9.18618851503935,
  10.2854237675064, 3.77193929847013, 1.77169185522596, 1.36923492824198, 
    -2.80974583059541, 0.578788004219774, 8.04495504253323, 8.86483075818995, 
    -0.60386414907931, 3.38714079495014, 3.808662360479, 1.15288002935914, 
    4.85007050264088, 9.44705845188831, 0.40486430955144, 0.303887155466496, 
    0.927426137236625, 0.041763927582279, 2.20267449810382, 6.9373296912485, 
    3.70846844704205, -4.35959339359339, -0.675214150407721, 
    -0.281611142284804, 8.82345218585665, 6.89799210505276, 
    -0.377106490829522, 2.29438354730976, -1.31713776609594, 1.0850637919515, 
    2.29661464418177, 4.67180436659448, 6.8305309707591, -0.87869263430519, 
    -1.55741293119148, 2.65302821447819,
  9.17011481490153, 0.600313473077633, -1.9664465213305, 0.21132646992456, 
    2.31278565550068, 7.84109727840372, 1.45780070877382, 0.188724145091831, 
    4.70349975541547, 6.48549368969597, -1.25763322092449, 5.5186866748489, 
    4.25571210146783, 2.00345011088195, 5.75040955294341, 0.214151038408601, 
    0.354304756783542, -0.672663513113145, 1.15229695996695, 
    8.31766817415136, 5.48492045683532, 3.06822327238277, 3.62807518696073, 
    -2.66563912817155, 2.55772088807105, 8.47804608887746, 5.75043321097507, 
    -0.0401773317866221, -0.17213165262954, -1.19641704530409, 
    1.67089444048029, 6.718820096361, 7.30025537166582, 0.0262751218307589, 
    -0.672914019101897, 3.56419506054874,
  4.5319912360154, 4.55155981538975, 8.91953839953641, 3.36433135575815, 
    0.799938234511923, 5.7626395970211, 0.0575925161343136, 
    -1.90223496412651, 0.507571634556503, 7.01318799636022, 
    0.385170762470356, -1.06762399041595, 1.04134725639591, 8.57025322474326, 
    -3.72918387431163, -1.20915720946376, 0.538402256035207, 
    3.77320854906553, 7.56077087532276, -1.42537177909716, 0.10585198125732, 
    2.21163257256874, 10.6024662977624, 0.856887957098285, 0.316768250846791, 
    2.39081041954518, 2.19054576582392, 4.34963090590086, 6.74524797464165, 
    -2.21927686775944, 0.891330451740912, 1.5920683646017, 4.82404243324885, 
    3.97499084987289, -3.81932239890775, 3.67521371083257,
  0.104962429844861, -2.12687586683223, 4.21360318102819, 6.71916385923067, 
    4.68584902468631, 7.16059776833712, 3.54600821199611, -2.58818539868935, 
    3.98221458822232, 2.48642701822042, 0.871351821479379, 2.52061306581946, 
    5.17567923438437, 4.97437595695513, -2.68797019071565, -1.96904342349394, 
    -0.547267231225241, 8.55623499480169, 7.2037952667645, -2.25714961924104, 
    1.54138222864364, 0.351048122236579, 1.18760470967471, 2.75244355403838, 
    5.8595338230394, 4.76205814098935, -2.63548895166815, 0.976087436569593, 
    4.15051703367317, 8.3550788433999, -1.72220945553321, 2.52402817158243, 
    0.937407668615843, 2.83945920034322, 7.14006087783144, 9.27779750529217,
  4.51202304309183, 7.93702366080283, -2.404757726133, 2.6956181680246, 
    0.227449338211951, 2.49946006255581, 9.64049118174085, 2.94979027444538, 
    -1.65319179795322, 1.96951561397708, 7.12947142709657, 6.42138275939877, 
    1.75882427948047, 5.58221724450885, 5.13450060538492, -0.130172982578008, 
    4.30219075244315, 5.42525097380703, 0.790939380435421, 4.90993687740627, 
    -0.227117876046365, 0.158427031518079, 7.09259282238211, 
    11.2427188927432, -1.81997141126422, 4.39142299031651, 8.03591574041772, 
    3.7569985548515, -0.883002513866972, 0.930012185177567, 5.35361178356489, 
    9.11348140099258, 2.33850692698084, 1.56238390723509, 1.229397658204, 
    0.846558657871926,
  7.39826236977752, 4.06638077121755, -1.9682309317159, 0.602627779875925, 
    2.92099084068737, 10.957396445024, 2.666597725926, 1.33821242411406, 
    7.10675681381474, 0.601620492499797, -4.47206305481751, 0.86996162570328, 
    4.23405488867767, 7.38095484842114, 4.91937202426499, 2.526813360845, 
    -0.0875716422579322, -3.39736705556332, 0.92628067432025, 
    8.28276281065279, 10.6849292635032, 1.91503962227107, 1.42433017228751, 
    2.8262292615284, -2.24620808801441, 1.90345003744676, 3.53609988445346, 
    7.80472076327119, -1.59128452955258, -4.04599698930156, 0.42219485667189, 
    8.28268270985716, 1.81849529510217, -2.61846405219182, -0.52722937334696, 
    2.38613521858918,
  6.21525949906128, 5.55957189593332, -3.5540253385264, 2.09936921441863, 
    0.200155325405332, 1.66380294800623, 7.19033709024881, 4.69398612562699, 
    -3.83737490784867, 0.0414990732165856, 2.55053151493694, 
    10.0703522589885, 3.84115912091071, 1.17972278881007, 2.25101178885747, 
    -2.58317341821406, 0.759151905130023, 2.18600096157601, 5.83467299307778, 
    8.6993676043306, 1.16474939522947, -0.102700828664698, 6.16853869618928, 
    3.77125335800048, -0.578416349788675, 2.54180582489901, 7.72651758333183, 
    -1.16527348741801, -0.293360932505388, 3.69220395697847, 10.016256512881, 
    1.85302519508958, 0.238510863950725, -1.29728904878637, 
    -0.492789233340532, -0.0696265325571388,
  1.70775984160729, 4.83774225889027, 8.16070125503315, -1.87189231382869, 
    1.13214073554666, 6.50439343115941, 3.78596825618709, -1.18150254039635, 
    4.57661096935633, 9.47935905703458, 2.85683694350229, 1.95393145927906, 
    -0.454969862871976, -1.93943636520782, -0.0441547711079746, 
    7.62974792367301, 4.78641783376311, -3.82708759684248, 1.81936360374852, 
    0.374297187708856, 1.77777513181007, 4.57195718788782, 6.04165766655469, 
    0.437360034582897, -2.81249690931, 0.77190053406563, 2.31243073491588, 
    7.88907305816462, 5.22928180011453, -3.33277525879157, 1.87820179922377, 
    9.11106757587618, 1.96367666550675, -2.47894605298626, 5.01296742877353, 
    6.16701280142242,
  -0.736999247281922, 1.34417159040163, 7.1233691385808, 7.43314144903977, 
    0.543153396082938, 4.38118767507898, 6.57968894788378, 
    -0.615931337051654, -0.65217353237193, -1.11675086336254, 
    0.822392075789724, 3.1051574870489, 7.41296821524022, 6.58639683278601, 
    -2.75512493608469, 0.929014943851669, 5.29262087512218, 2.7725366809325, 
    -1.18167985498248, 2.44811835522022, 7.45094869607591, 
    -0.905806067616421, -1.28764858619468, 1.65558279213732, 
    5.74211342547532, 3.38682360418955, -3.32972058964697, 1.06996384596986, 
    1.75497514102092, 5.84003063377281, 4.28954731864197, -3.00870170762094, 
    0.749808144862593, 2.69734094419296, 8.00250764251094, -1.2405684981108,
  -1.90841925406193, 0.719787376758258, 1.53160256100566, 5.14477963445267, 
    3.56820163376692, -2.96645397544719, 3.40749509084772, 6.66576595580935, 
    5.04305321664825, -0.351885474041083, -4.33722385229735, 
    2.16620748689413, 2.0248535926747, 5.12789631281529, 9.48164804264288, 
    0.456748080186162, 3.04605775263318, 3.26888751957784, 1.19623842295078, 
    3.9511847349346, 6.94887462038904, -2.91196533262478, 0.278093479547418, 
    2.18618899056182, 10.03940871384, -0.526458175066058, -3.51877093084022, 
    -0.680864261034496, 1.54769264978549, 9.1264925306793, 2.93999208978048, 
    -2.03732187080591, 0.420460971808732, 0.802297792003434, 
    3.23982738041944, 8.33686259558307,
  3.54804396476376, 8.30063907959056, -0.784158280312655, -2.63761947699717, 
    -0.0840662445803182, 7.92282242954595, 3.91393194490572, 
    -3.61777676849146, 4.05593368824496, 6.10510031342412, 4.40502689332365, 
    4.43550900912886, -2.21967310360057, -3.21107572719003, 1.76779157388924, 
    3.91919312476553, 3.29404415668741, 7.38766042148701, 2.6153010213113, 
    -1.76189211193214, 5.34215677947124, 7.84512014579138, 3.46913997415469, 
    3.25485243367415, -2.47708134393021, -2.01157540772967, 
    0.433799279991173, 5.32384618767109, 5.33559460725486, -3.49598302560114, 
    0.305702083180657, 1.1832643341122, 4.59452849485344, 5.41332312420785, 
    -2.65440445850268, 2.18209432065365,
  0.173199145194658, -2.64669323933657, 2.11249850231618, 6.59608723599963, 
    6.13878183894822, 2.85319039686404, 0.0361748468081839, 
    -0.390404046113666, 4.025848438417, 10.5001475514672, 2.81146897599318, 
    1.63279003904593, 4.32602171840234, 1.88562479863403, -1.25082110339009, 
    0.701578521708696, 1.64090789760614, 7.64493121589593, -1.71074738177969, 
    -2.66306938794912, 1.29326550729911, 3.90502622871383, 6.36400552273382, 
    7.35930101688194, -1.39950625027323, -0.661050730189674, 
    2.13946018488786, 2.23447683641469, 3.50850435582319, 6.13055021503629, 
    -2.12513910259206, -4.07272069353652, 0.162928502144271, 
    6.06429532228625, 7.02139167060585, 4.01300507353037,
  8.60591013077017, -4.67972804708293, 3.15401175916151, -0.449675007748443, 
    6.05734079464004, 7.39522661689649, 0.56478248881394, 4.72526066489942, 
    0.589177615367722, -1.11514936768, 1.05375810035858, 7.85906452178346, 
    0.596264220868541, -5.22324457235125, 1.03103416946575, 3.23054610738313, 
    6.84588046108741, 1.73828450195548, -2.51565985790279, 0.465826781154799, 
    2.15081117480586, 7.8179482978515, -1.02955484506679, -2.31645404707626, 
    0.811407250683604, 2.85886225623211, 5.81872451358078, 2.57229914015316, 
    -3.45718490906073, 0.860910715454938, 1.42429161628635, 8.67835622184662, 
    0.701345444076067, -2.48742488077634, 0.754880510846866, 3.44352817142283,
  1.38116002246341, 7.47096680772888, -1.41062197665313, 0.244302328325435, 
    -0.837269723548457, 5.97425645292102, 7.27611772054782, 
    -2.53946086954017, 3.01902957861591, 3.22288354164254, 5.37025805659041, 
    6.21132519230183, -3.88263920533404, 2.96696493672938, 4.44468014512288, 
    8.08140879893469, 0.34298526546732, 1.89683912143914, 7.19989583048246, 
    10.153020982481, 2.33573922983588, 3.63423823780623, 2.41735887010706, 
    -1.69745343871194, 3.0630091857896, 5.25274283332612, 5.97712760206098, 
    4.47888318216297, -1.03103984819697, 2.91203987300318, 9.5710676614072, 
    -0.967541125813891, -1.59276001204821, 4.75804556788352, 
    4.00269834952864, 0.0867382896723634,
  -0.941300593054871, -1.21240559206636, -0.256248493878743, 
    9.67948421145043, 8.81086042019873, 2.3011313171475, 6.16236073227066, 
    -1.29745220912424, -0.248420764406888, 4.32519709696589, 
    4.47066842374646, -1.65921503136642, 2.12556034215197, 8.29659131727636, 
    -0.293330731994694, -2.90997601888021, 0.813755284059162, 
    10.1989027728437, 0.549380680313609, -4.32569975345797, 
    -0.0613324654355751, 5.7158471867142, 4.5477842784643, 0.31009743030107, 
    4.27583387595321, 6.37364946820163, -1.66627844927751, 3.51917597639907, 
    3.4167756473824, 3.70475203359751, 5.62626044484867, -2.58042943339981, 
    -2.91832494771653, 1.42560604369949, 5.29477290480467, 5.33827420841603,
  -5.48659823040787, 2.37431907641058, 0.238425853254594, 2.95820000845448, 
    9.28393428881868, -1.91428516939276, -0.0997966767850076, 
    0.817430814891702, 3.38188962776196, 9.425369358943, -1.0689950396786, 
    -2.41957450401426, 3.81695066182224, 5.57242368610171, 0.417359016307493, 
    3.50422201354255, 8.44853190083081, -3.01328628762143, 0.301185515039166, 
    0.582222105898422, 5.64883430492051, 5.19845920654572, -3.09400378155233, 
    4.32844339166365, 5.09572989741311, 5.56103521262436, 7.07424032034198, 
    -2.09854714368814, 3.15061708183273, 3.84422416368865, 5.33418324409706, 
    6.95672180728995, 0.776678355235165, -0.137340286753876, 
    4.38400597235317, 5.3830962006534,
  3.21229312004672, 8.80900846518104, -3.17598801490038, 1.45865018812989, 
    -0.0663389646538874, 6.1150105615109, 1.11988819763428, 
    -3.24117286537152, -1.64486474956226, 7.79283717458398, 2.48674122071749, 
    0.217037285506516, 3.14059512755109, 10.9370890292885, 
    -0.466235912781947, 1.3211940046189, 3.80997513607933, 4.94426843211768, 
    4.68972130369503, 1.511094953267, -1.1848952123696, 3.1096675756015, 
    8.65126829905972, -0.263158939123628, -1.93105803580787, 
    -0.766564824031992, 1.33144798079557, 7.19968613307704, 5.37815291670085, 
    -4.47866095964547, 2.64808990924387, 5.89407693194526, 7.10512997056657, 
    -0.10650741337214, -2.28358122831848, 0.0656293759217257,
  -2.26053384657504, -1.39894356477956, 1.2172009786682, 3.61667165663095, 
    5.578051838303, 2.63462181569816, -2.52727776197206, 2.05295175832984, 
    4.32147567494906, 5.79364807867712, -2.32877327090298, -1.69187927481553, 
    0.561864168867597, 5.16208220576554, 6.89661610868855, -1.91717272540117, 
    -1.83532460322114, 0.411855220939949, 1.55013681191917, 3.82528592648332, 
    6.13713528037427, -2.08431243883018, -1.62384484145975, 
    0.573477106034121, 6.55619123746178, 6.80313460898412, -2.90320531976946, 
    3.44840053615789, 5.95652208972871, 4.97445259867809, 3.7750736706356, 
    0.525523402276585, -2.02816968658542, 1.82671689920697, 5.13258847973834, 
    6.56189683753603,
  -2.42534230300052, 4.06814729951094, 7.37698943655106, 3.78385926780482, 
    1.55683847048705, -3.12498112945861, 2.40846291187213, 1.68737622051058, 
    6.11556678735472, 3.85260305007899, -0.809539547189326, 3.57803153578832, 
    7.78566356587456, 0.390059846063603, 4.31923688011655, 7.64889269255612, 
    5.15773862834554, 0.908288006682996, -2.03609683075925, 1.17792779629832, 
    6.44294531473483, 5.80874538972708, -2.36131224868884, 4.80917840120181, 
    3.77371729138971, 2.64322380353972, 5.03061271026087, 3.52072585159471, 
    -3.1139843744322, 2.17444934032104, 1.51919770346328, 7.1390422564288, 
    7.66875471057068, -0.593124285568955, 6.27754069828341, 4.38283829825322,
  3.7046595041378, 2.68142789903841, 2.66641142853334, 0.0677340295031845, 
    -0.840627408700016, 2.48658019793757, 5.94774262736231, 5.7341423157767, 
    4.58473737971601, -1.24724042720268, 0.559529876802864, 3.4138834844922, 
    11.7669658159759, 0.805925725159402, 1.24466411320473, 5.09333208841553, 
    1.82052325163404, 3.21941846806765, 6.79359394224319, 1.32511670884429, 
    -1.08575372120692, 3.09387743402114, 8.96610308440844, -2.40996287639269, 
    -0.76523017162508, -0.269428813584268, 0.477109295296905, 
    0.911236176242876, 7.95078714376618, -1.61621708998508, 
    -3.55709160221816, -0.68399982353098, 4.59503591699917, 12.5983371222375, 
    5.58056656690628, 0.376622597535755,
  -0.911687177642509, 5.16836849631074, 8.66682364032584, 3.44948207502787, 
    1.72656668319968, -0.923102964900454, 1.03193669316399, 4.06334641735249, 
    6.63354864126004, -1.79412806913545, 3.48457520160496, 7.19262737270035, 
    5.18711633357535, -3.098116331708, 3.92130032943168, 4.56550210909592, 
    6.21289964429401, 2.4297013446692, -1.08497357257359, 2.7227405659925, 
    11.1559755029662, 1.13424531884868, 2.98446754524002, 6.00223799959071, 
    -3.49466163102194, 0.377443580906831, 0.519913516559707, 
    6.19561622213323, 8.58562105654171, 1.38923147938815, 0.377953751830777, 
    -0.106452269654878, 0.155435161545013, 1.70566828314297, 
    7.94008644722685, 5.65392722475764,
  4.4212273444717, -1.48837431220816, -2.75324354146435, 1.16462772952946, 
    3.58141965887477, 7.38108412495674, -1.36051995419247, -2.79030098116668, 
    0.667483811799845, 4.03158751505027, 7.00518722896905, -2.54925808048095, 
    -0.0633588755782295, 0.530841937347698, 10.1757025903346, 
    1.0239018616751, -1.36763497388101, 3.80351649092544, 6.27131937303085, 
    -2.87172890005357, 3.21246371541414, 3.43843110565666, 4.31185918147784, 
    7.7236375516002, 2.4745220369793, -1.03812572811969, 4.46991809726978, 
    6.52864212779784, -3.10523834922317, 2.17133575523527, 2.29232230928413, 
    3.83112241815835, 6.8206057606306, 0.169092851266708, 3.17731686353642, 
    5.36296296423816,
  6.6876532615221, 1.86622426773716, 5.74003662223128, 4.8859714210637, 
    -3.37507342917583, 0.246494431568369, 0.70961153668621, 2.41955496581664, 
    5.48370991726688, 4.29935258857824, -2.86564549605245, 0.441739301119287, 
    1.66277386668616, 9.03632910589625, -2.04085533759722, -1.69846341075455, 
    -0.613128984357575, 3.80728294756364, 11.1565283676713, 
    0.587148420182069, 1.12235243949258, 1.78091790165564, 0.658636281325161, 
    4.06456948206796, 7.89053934097411, 4.08803704215639, 3.22317700191125, 
    1.57646696322298, -2.20214791614842, 2.25842772789975, 5.82627112938011, 
    4.56201527978935, -4.47563333925449, 1.36326380425524, -2.28270450056296, 
    7.14351225281251,
  -1.38598499125038, 0.441848927520351, 7.25756691811712, 4.43242251162876, 
    -2.73784755290306, -0.623735910974469, 1.56743896036054, 9.1238488534374, 
    4.29226776307009, -5.70602359399999, 1.38395588576834, 7.02890175538225, 
    5.89548947656166, -3.46871611745881, 2.21453768684672, 6.54567167346465, 
    0.79150455823221, -4.28206088638595, 0.378672209986414, 8.67739225000739, 
    5.31701263244431, 0.532852248992407, 4.96614704595793, 3.24404662118201, 
    -2.16831726823503, 3.77449092850701, 3.80649473217422, 3.30633096049039, 
    5.9098205244512, 1.94869386433028, -2.81129987605936, -0.412974641650192, 
    1.94533492612131, 6.94091785108462, 2.6181494779659, -2.87098545693273,
  1.87603550851618, -1.01742605545171, 3.55572008426513, 8.63630352073437, 
    -2.92301232166407, -0.570702250669516, -0.527738919314352, 
    1.00777445627867, 3.23824162475187, 7.2890678454548, 4.20663810953409, 
    -3.43106285882501, 3.33914601243268, 7.10067922240326, 4.19300924001698, 
    4.555406683053, 4.05041643114706, -3.11893106084497, 0.459069021342257, 
    1.107518452843, 5.46485792228791, 5.14513350546994, -6.05329001699045, 
    1.05243732552328, 0.0983568901142191, -0.170684594075419, 
    2.79479009855731, 8.65305681334815, 1.04838636124126, 3.57135214652502, 
    7.07315521513502, 2.99688142858156, -2.08629815322078, 
    -0.434755368033996, 1.67645857179334, 7.83846709550656,
  -2.50902161162322, 0.309615073589232, 1.856825170185, 9.01896691212908, 
    -1.6926651675152, 1.59408411928854, 0.721072061124896, 2.16114021377106, 
    9.26065940386391, -3.76563923382541, -1.3296140404736, 
    -0.626681641679208, 2.71799698123904, 9.24512296086119, 4.93774410026696, 
    2.32266699621456, 3.48655891075609, -2.0640600851905, 0.480473703660265, 
    1.30393888916366, 3.36785923849102, 6.81431566562649, -0.340130741418215, 
    -0.950574376945099, 2.55621073089117, 11.9807237445141, 4.02860172228928, 
    -1.18291877059965, 1.72267353568003, 0.541512786064537, 3.61058799497477, 
    6.23877895925293, -0.952496684330314, 2.52173692631881, 5.18134881631081, 
    5.8978997099901,
  -2.18469765989102, 2.87040292950078, 3.72727192462834, 4.83686944127653, 
    3.94183459498183, -4.21236792347453, 2.7682864110067, 3.12578303472749, 
    4.23061010046316, 6.52479812866186, 1.36335589132683, -4.44436465013949, 
    1.60777868177225, 4.68301566774025, 6.1017859880767, 5.39566648201831, 
    0.252687658513727, -4.1526797973705, 1.70633341923743, 3.75778639859217, 
    4.7556912487063, 6.53834737792508, 3.90745912808882, -3.19136793993095, 
    -1.2812347141252, -0.305641658379173, 1.07581851453777, 1.83998048895525, 
    6.04462838469141, 8.74758436879626, -0.367963324215212, 3.43975389888139, 
    3.36944410187277, 1.85711015090987, 4.31002129856333, 5.34714800471795,
  3.06958407304734, 5.76539962800815, 4.50306635651055, 3.98576847199181, 
    1.32421821015954, -2.93771674639315, 2.39948790896968, 4.49240031926584, 
    6.53716942090894, -1.90746763636172, -3.77565056662208, 
    -0.84003567265814, 9.07053645364011, 6.53510679717011, 0.992295493047792, 
    2.08572320020153, -1.5504367726121, 1.76561123361767, 4.4726819476746, 
    8.86490552607349, 3.65636194216489, -1.19888881922078, 4.93325091618436, 
    7.92752118714758, -2.35199655932499, 1.75217318019771, 1.26162451004547, 
    3.21633248255447, 9.21116131271996, 4.7444433058349, -2.34242959787116, 
    3.72293755602125, 10.1406183071962, -0.896757155635137, 
    -2.76027907445774, 0.367795588017065,
  4.76446950029741, 3.45763068531338, -1.72194937763132, -1.38066531536416, 
    1.07056850616769, 5.35166901983091, 6.29139387607121, -3.72662328824996, 
    -1.92823263755439, -1.67081659546407, 6.89873669442963, 
    0.837348185855494, -0.736455687269031, -0.332562040325391, 
    9.64965100396761, 1.29041295510428, 0.686262951551335, 0.895047112381717, 
    1.63006887625475, 6.88607453692175, 2.62244420497603, -3.90962567761403, 
    3.86934124093055, 3.78734919843657, 3.32219669377162, 8.0436899569226, 
    -2.77982621137225, -0.166894231290359, 2.17587254354308, 
    6.97250901248229, 5.37520076417358, 3.72056581507026, 1.27841073652487, 
    -1.70199771578773, 3.10857751540068, 5.6171058513049,
  0.834689881547722, -1.06368893038716, 1.38687156495146, 8.98649991960819, 
    2.28059034978829, -3.9771586911168, 0.268030571520379, 
    0.0422584577913168, 0.372400037260379, 8.33576248376454, 4.8457516381552, 
    -3.45305903684207, 4.30733633162866, 2.51112369123641, 2.39755650772127, 
    4.95503953611581, 6.23354641820551, -2.16765213367698, 0.141017850778114, 
    3.52226524772148, 11.9927552122202, 5.03444337829477, 1.48068765023908, 
    3.40443452634891, -0.93110799474572, 1.85939310159392, 9.60002467508417, 
    1.88453578967746, -2.33965694206259, 4.02173011261262, 11.4807634614671, 
    4.01708114030035, 2.90599298514945, 2.95008104194761, 1.65353760806642, 
    4.84663651133838,
  -1.40267161236462, 0.790129465913728, 5.24058683144902, 2.62069056971511, 
    -2.39626130073295, 2.10125378284434, 8.35626317749679, 
    -0.154504009781772, -2.47356372688727, 0.713562892289822, 
    2.58133301078728, 6.5225541126488, 0.493816281019705, -3.6922625926326, 
    2.65269172869787, 10.0899212643419, 5.00387962745714, 0.197086578435461, 
    1.54963720372876, 5.64442290226905, 2.15813304544779, -2.50705298860919, 
    2.93713285867772, 6.19425227960742, 5.62194660007359, 2.14532163487786, 
    -4.00265397550307, 3.10443665434396, 4.21710276774813, 5.3093812105629, 
    0.894297039160687, -2.68282025776847, 2.58222714999539, 7.11170941438876, 
    6.41856823245402, 3.67450004051328,
  7.63024291656427, 4.58470837588697, -4.46149971288154, 0.431285364795389, 
    1.90450660764772, 2.80362758306415, 4.07719293229708, 6.10350435468817, 
    -0.669107693963445, -1.33769282621349, 2.23134807210681, 
    9.49481399750958, 2.79367217900059, -1.75128421103595, -0.77023169597213, 
    -0.13236673071459, 1.42984398358757, 5.52895317140468, 5.80456995041007, 
    -3.26202901350711, 0.991841062766437, 3.96650526766873, 6.44391698922401, 
    -0.304644349981328, 4.86267416546601, 10.3270022794557, 4.97701378114051, 
    -0.519793007134451, -1.33691394744198, 3.55792105587248, 
    6.94576730323295, 3.40219169862269, 3.94913181382282, 2.48665836005266, 
    -2.17991090759827, 2.24980711781576,
  -1.84426740050893, 1.59723898793408, 0.688299425181985, 2.78474920940806, 
    6.59910459344163, 0.865224904420662, -2.35276304081077, 2.67943362935658, 
    7.02182141227337, 3.16979324798564, -3.7448221910451, 0.993755152797004, 
    -0.0103928441710872, 6.98523551174885, 6.62174080815964, 
    0.0134807171220528, 5.53561209803696, 0.784789952222282, 
    -1.2129674933411, 1.062274151727, 9.46100217395366, 0.503532404817185, 
    -2.17032210732846, -0.792788937019142, 1.42817104591156, 
    4.85699188951688, 5.8727662677719, 0.268478238250955, -2.09040282300205, 
    2.4854065354679, 7.366142469106, 5.88393913972516, -0.656775864968888, 
    -0.211122151592708, 4.40466319189974, 9.04114984200016,
  1.66041065962136, 5.99708771562321, 2.91046829588175, 2.82217479408147, 
    5.71614174315929, 2.682521933812, -1.2625646362949, 2.96603761505432, 
    7.54511158973639, -0.324233051700091, -2.98323223547867, 
    1.23456978599996, 2.41805748104784, 4.55366569724953, 5.6879077676338, 
    -2.52424562106928, 2.75094998700851, 3.06368151620952, 5.61184942650907, 
    6.28855675713334, -0.890521610363816, 4.25691707887589, 6.12731446153427, 
    4.54971387701256, 2.59185973018471, -2.01360800970488, 0.995492635487021, 
    2.79389381867085, 6.17375454341569, -4.11505195220321, 1.03161234408709, 
    0.622294568519544, 5.24123787936708, 9.45478047887592, 
    0.00352295229310862, -3.17539621051294,
  1.43328300430001, 7.3794106718332, 9.01867093792166, -0.116334321641274, 
    5.65775401382775, 2.03651036981519, -3.4431355793675, 1.22984170210519, 
    4.42510259425796, 5.64533641639122, 4.2491664706004, 1.15717787175934, 
    -2.69268876081461, -0.316333859008319, 1.79199251615802, 
    8.94524271470391, 4.80532340823676, -3.23827571199136, 1.00265692911026, 
    5.77928433398557, 1.04069667897932, -2.53972666704467, 2.07249508465085, 
    7.86102138739943, 7.20540001582631, 2.71218392994724, -0.691943816885837, 
    2.78451935987093, 6.57870142360813, -0.874415162522492, 
    -2.45697316789154, 1.73943774921396, 6.05057364559897, 4.63181252178881, 
    -1.72481586766041, 1.5825121455922,
  2.94295132859482, 4.85046837563234, 4.35765244827041, -2.73211749362781, 
    1.89417884864578, 2.66384269199877, 7.50178362920831, 1.86853258328623, 
    -1.73008306912009, 3.32301514290059, 8.63871429502431, 
    -0.662230100938016, -0.557094507868849, -0.790018547765216, 
    1.50300140413202, 7.36349635459242, 4.09829072631755, -3.38271512342639, 
    -1.08345910887143, 0.863889394776344, 2.17256848132286, 4.02111481072152, 
    6.77720305642728, -3.30460725005257, -1.96464497487748, 
    -2.33946655516074, 9.13533360101896, -0.116498718280043, 
    -1.15173667706535, 1.52158561552711, 3.42204268501782, 6.09399347229029, 
    5.72276565982372, -3.35022147476214, 1.69949323028902, 2.20640502469513,
  1.22210066263062, 7.64979116588753, 6.29450207625883, -2.55301058955779, 
    1.03363288550253, 5.66176651106371, 3.16853325106798, -2.83401476101341, 
    3.58526560694988, 6.01098532452038, 5.54570884009392, 4.13017920047844, 
    -3.04827459850637, 1.34278924482342, 1.12458121403411, 2.52797679779249, 
    5.94460253725179, 2.67407601378663, -3.51764252481681, 1.42802550639049, 
    2.13740875298609, 4.87547574033157, 4.99492251343351, -4.00941976116042, 
    0.892490004190128, 1.59196597858598, 4.63567495387325, 6.28938339445215, 
    2.64718013929137, -1.68844686102749, -0.42441032136047, 1.86182688293503, 
    6.07382014199944, 3.94961515294312, -2.63253177899101, -0.549515683318476,
  0.538472186184307, 1.71910658333921, 5.28907628959396, 6.16801415008183, 
    -1.81813432238379, 3.8188053786305, 5.36817749584585, 5.58036372759192, 
    4.76469597074176, -2.71314628840778, 1.1299910196964, 4.37067005131208, 
    10.0706814970518, -1.28257045370596, 2.71722468225248, 2.6805011610408, 
    2.02521042771675, 3.65652698580662, 6.05292989460368, 1.24033157425983, 
    -2.64527082601309, 0.783967751773949, 2.35977964448635, 6.42712976537664, 
    1.215586554244, -3.91475094958942, 1.30671162098142, 2.7150866674369, 
    6.80848483270399, 2.35745470501945, -3.91403743144087, 0.764770800882509, 
    2.70663730957273, 8.75683916713526, 0.517873468418449, -2.48930273398165,
  4.96275292837505, 4.89771792255423, -3.05843241422803, 2.75454461221682, 
    1.98566334523829, 2.92703894104953, 6.40282655564083, -0.334267231769557, 
    -2.5578201970606, 0.912045088760461, 3.58160135377335, 9.22164507764056, 
    -3.17237976395229, -2.08296267228015, -0.870105206198208, 
    6.41114229697392, 5.43506067717638, 0.594210777010576, 4.62776943388108, 
    2.85576546983855, -1.97335334554873, 2.90589161905659, 6.87034721097885, 
    4.1093078572822, -0.0890866480197095, -2.20402911831801, 
    1.35651031393112, 3.51712162261671, 7.10739939155223, 1.80090205826706, 
    -4.04583257131427, 0.853905220487193, 1.37358731852407, 5.98924221722807, 
    7.08005806144525, 1.52562570733193,
  3.31894350302585, 9.08772217527211, 2.67493116519076, -0.411435255227798, 
    1.11263116335626, 0.519167061534442, 2.63619824075016, 7.26311057079933, 
    -1.37264902362671, -1.51844512211675, 0.887565436827336, 
    4.19321403747136, 6.30635536626483, -2.51721459593611, -0.36585337312354, 
    1.02176967906828, 5.3873922722425, 6.37044513745385, -1.68317291868729, 
    3.70724975387223, 4.93205942272596, 5.26127487330336, 3.86711471959822, 
    -3.04018217361767, 3.15893365716225, 4.49904358662273, 5.45617242225213, 
    5.09170900720063, -2.57495555856743, 0.566110900154893, 4.35241298741465, 
    11.0631558010435, 0.253113229474585, 1.00869552217871, 0.955926005370138, 
    0.456137386792763,
  -0.270647613159146, -3.15881988746445, 3.04095008510035, 2.18370212665153, 
    1.8065843232806, 6.62963685971598, 1.09170883874225, -3.33931082014541, 
    1.36079278373737, 7.02898233160652, 8.19481570099273, 0.28315929273302, 
    3.55882465515021, 5.24482397914896, 4.33930905860698, 4.99557699451323, 
    3.21095496717488, -0.0149571964264452, 3.62058704047767, 
    7.43171523320079, 0.200377092232013, -2.7862177021015, 
    -0.042225640644979, 1.35555546678667, 3.98761461241555, 6.52933496314947, 
    -1.18757591915257, -2.089164598411, 1.93327702250258, 7.57326567132888, 
    3.79636218604424, -1.39308873381735, -2.08930380691824, 1.66252882536082, 
    4.67540366562198, 5.87315475389931,
  6.92646389957976, -1.6789603137201, -1.82827297238235, 2.1686535050811, 
    4.09929126759172, 4.7453549170441, 3.74934536591981, -3.18564461888381, 
    0.80585803793664, 0.998913914109495, 3.19320695194786, 7.76995051629983, 
    -0.439852776710199, -4.11359787758539, 0.124226681233789, 
    5.5666008490275, 8.60033595330775, 1.66142595882453, 2.40232438839732, 
    1.23342536583329, -1.49791793586591, 1.58412518902075, 5.24081899139288, 
    5.55426586452225, -2.62958365466391, -0.180478853171552, 
    1.09333457808166, 8.66956340146371, 2.86592338559314, -6.26325894308442, 
    1.08498657191956, 6.66665543816473, 1.4941252388357, -3.51815413396291, 
    1.87451219574041, 5.24568115496921,
  -0.843833242314221, 4.97878552098806, 6.01003470025122, -0.368699331265794, 
    3.94946303337491, 5.95894007070532, -2.15427930825691, 3.51692291373534, 
    3.90207959910647, 3.9615882500387, 5.02312906913269, -2.31652149750434, 
    -1.25925665108482, 0.961394397128366, 7.9702395043913, 7.66098353855348, 
    -1.87438052393877, 1.8305148642245, 8.00123857295522, 4.86607094621467, 
    -1.00661848672154, 5.81665508502766, 2.42191335670157, -1.41663634338662, 
    2.11763799468147, 8.93203036907766, 8.49245517113436, 0.190132299804894, 
    -0.936262541171696, -0.348338633232996, 4.00368813527111, 
    3.47261734711111, -0.304703477833102, 1.57617880875117, 9.04302101392591, 
    0.24458138526692,
  6.6977480179396, 0.773202838401269, 2.43403335248495, 5.69477057662795, 
    9.96254776253402, 1.47777618845191, 1.65336292219464, 6.16763662908019, 
    0.360234827458124, -2.46126830353711, 1.06804529844322, 1.41411718321376, 
    4.575949208627, 7.72421555388567, -3.46380967652177, 1.93851250400681, 
    0.142415187209908, 1.68489656639363, 0.796838370094469, 3.00149548661285, 
    12.2195630959223, 5.028962819096, 1.85184745670326, 6.62971322462887, 
    6.70458618391374, 3.90938645653379, 0.99381418219925, 1.27128930354099, 
    5.51460735322799, 1.6758229051675, -1.20748462218903, 0.594643367484046, 
    11.6304930246522, -1.97368857936625, 1.08378066614799, 1.99590452987782,
  0.936514006605796, 1.56919583107175, 5.38854729488728, 6.56891869006337, 
    -0.340635277585441, 4.97008367191881, 5.77508985537804, 4.67555403418803, 
    5.52282252176533, -3.01244657911011, -0.30345286354339, 1.81576619869926, 
    6.57369701313936, 4.60625417774878, -1.88134281834534, -1.57803972405257, 
    1.98810994240621, 8.50430941011765, 6.80964993771987, 0.551665098966232, 
    -1.50504268604978, 2.55539455282152, 7.85995944461722, 5.00482011143216, 
    -1.45647012990436, -0.154755417301922, 0.574386993177161, 
    3.3483681150384, 7.53864694932818, -1.55981342181168, -1.43179196428067, 
    0.0829888202581426, 1.96673657680639, 8.43125004113949, 1.47421380694337, 
    -4.24409679920361,
  7.30232865021503, -0.507482914253751, -3.34152214905366, 
    -0.707394466831346, 9.80414036207154, 3.55015827613669, 
    -2.48636833927625, 0.851121365604552, 3.66557677791271, 10.3035715510592, 
    0.688982891398146, -2.2695783136201, 4.10653393674183, 6.31346314633913, 
    -0.853243534807207, 2.98311207232457, 3.36168289261988, 4.87040770602831, 
    8.1246838070533, 1.27493019635734, -3.65281158090286, 0.68600388425002, 
    6.94596999888484, 2.11973555535577, -1.45682363513227, 2.4415282455981, 
    9.2459081754301, -1.58644214853531, 1.86426536220382, 1.76239015778103, 
    4.38012552200903, 5.68194122007729, -4.4908428496146, 1.94496071625575, 
    2.25019426752627, 1.65906306270447,
  5.44515346596557, 3.6459734940711, -2.59003216116367, -0.995306339510443, 
    0.764968048123577, 8.11940696578688, 5.16725747415532, -2.94298517091133, 
    -0.0650016104938884, 1.22818469702442, 7.12397091153027, 
    4.36696943968822, -2.69467389103479, 4.23434186808605, 5.60626848542616, 
    4.14990598387873, 4.90644492464063, 0.179310157785587, -1.70736782284464, 
    2.37668919251938, 8.57777195265902, 6.32561459943124, 0.0913549948737726, 
    1.13862163920871, 5.83500431301939, 7.34999065740899, -0.142600527807458, 
    1.14842189943289, -0.263373369180318, 1.37341204965302, 2.91424834431913, 
    7.38864798558876, -1.87929475034875, -1.82773534254448, 1.40310284284831, 
    4.49475926472558,
  3.34020800902242, 5.12434710941299, 3.72926056457156, -2.66814047026142, 
    1.04484712180495, 2.30468212305106, 6.30884447355898, 0.817766111472072, 
    -3.51755588056716, 2.01566263625436, 3.97906661424346, 5.99089759105639, 
    5.90044442981691, -2.39848047868054, 0.159052902227519, 3.13904992146805, 
    10.255051990638, -0.64353486472661, -0.101283460017462, 1.77814860224845, 
    3.39700189160476, 6.71886577024239, 3.01902106466133, -3.85176700072843, 
    4.32825559172561, 3.84177924390028, 3.38812599873861, 7.99787560533131, 
    -1.52009270547554, -1.71583226021528, 1.93816748782919, 3.86605497484485, 
    5.04906091030495, 4.39663494693317, -2.5381567672479, 2.37650624719053,
  2.58290986283048, 2.25382587581638, 0.839083192374695, 2.53783823160693, 
    9.74880031709323, -3.92098053498703, -1.37865452433379, 
    -1.65472596984837, 7.07646963076039, 2.5683922457828, 0.554765618585238, 
    3.27050470261011, 10.6623843886073, 1.78047177187971, -0.55688207040782, 
    5.26110047864595, -0.745509836237526, 1.05272786083448, 1.53427899652402, 
    5.9682939335069, 6.38817209475325, -2.86210998894445, -0.227825356765015, 
    0.960881659874233, 9.83123013391498, 4.35417329269104, -2.60526396716791, 
    5.15860532758792, 6.87798283747445, -3.38347201174481, 4.31611333480607, 
    2.78029652853606, 2.00067420879908, 6.30074932391102, 7.61620047988331, 
    -2.60178435102468,
  7.3929872354349, 3.35674531856772, -1.44899444675094, -1.66807375057726, 
    0.947110935788993, 3.63646091916056, 7.91908474048545, -1.89171400871003, 
    -1.49698202246254, 0.542427484960889, 4.17965624850561, 8.23338645641395, 
    -1.76538866905099, -1.62786660178079, 0.426365468107942, 
    8.94707051205267, 3.77311201749002, 0.234133068468906, 6.12310318692115, 
    4.78531866295301, -1.630585769443, 4.8876452531355, 6.66405777887479, 
    3.91582165821452, 4.7275122184348, -1.27520334926072, -4.06511257857112, 
    1.94770940979486, 5.64466944650743, 6.54671491104577, 1.72078006523975, 
    0.0968357388165289, 4.56846467603879, 4.63900442743168, 
    -1.62147437231316, 3.3430096885105,
  1.36305144977287, 4.27899752349592, 5.54359723913362, -0.621590325091284, 
    -3.01949637362591, 1.34822488446723, 3.01050282358178, 5.51996111310345, 
    5.11210300935914, -2.63241450881387, 0.869204263238422, 2.30680384576127, 
    8.57086821223718, -2.3292093282444, 0.244829156714073, 0.542803261541956, 
    8.23634145270357, -1.52025146934061, -0.212001242578582, 
    0.904661012834906, 4.08998135702736, 7.69550041152081, -2.3354616463731, 
    3.46824274138604, 3.17402605507561, 3.44272293885773, 6.6453222581955, 
    4.29675111886849, -3.52009743432874, 3.0387500674784, 6.7234811375448, 
    5.04947244278689, 4.27107938634622, 2.69220985528344, -2.37378695844497, 
    -0.102241187261861,
  -3.69328330055333, 2.07132465072628, 6.23905079704422, 5.21121477550795, 
    -2.54205328635992, 2.16920823157081, 10.9153521090772, 1.11054562561237, 
    -1.44474597643087, 5.56990073231704, 2.43011360759196, -3.52881146136116, 
    -1.46781422614516, 9.36850226216174, 0.430011781719317, 
    0.677971395922222, 4.06298967412749, 6.06797144791255, 0.371119538852751, 
    3.29790292436483, 7.30595630903445, -0.364361700491831, 4.19060036411199, 
    7.03203174716697, 5.90054085663887, 4.15957586803393, 1.61047618116372, 
    -1.06869148392352, -1.66197382938528, 1.60479997555719, 4.54545623442041, 
    7.79046226160531, 1.24675803042373, 0.656128196763602, 4.79588197026609, 
    7.9909860828624,
  3.35582801330418, 6.96771116150938, 5.44193891176839, 2.640161864673, 
    0.144919876298858, -0.214991381515507, 3.40566293846176, 
    10.5949413049301, 1.77083612721471, -1.17903163073996, 1.51354910732762, 
    5.19390480486378, 3.95074151719148, -4.04047481018726, 2.04403378875775, 
    2.67748630557154, 7.18735186487428, -1.05458951578824, -2.84205528399086, 
    -1.33276606496148, 0.897520318127111, 6.31715827864272, 7.27839704674977, 
    1.44864105098428, 1.16183873573873, 5.38203426946378, 6.23337180322255, 
    1.56709526736547, 5.25842649572, 5.68619091360793, -4.47309645058485, 
    2.17637051417481, 1.58325546685778, 5.3138004657986, 10.5598464005846, 
    -0.74320424513781,
  -1.82264900722812, 0.158870919747497, 4.13635265668157, 6.36704303986705, 
    -0.00659553743261121, 1.81240446742124, 3.86970802512766, 
    6.12179878648323, -1.48262199138992, 1.97236565418944, 2.58376623580763, 
    5.79342408125806, 2.02564563821608, -2.26056981213639, 3.20935798801204, 
    9.14742820161201, 7.18118856176842, 3.75458092222904, 0.970984164556466, 
    2.75757787642538, 4.07383894061163, -1.28413167291236, 0.689586656633972, 
    2.02057298457301, 6.74327866222399, 5.56186486378852, -2.55640062209585, 
    0.283262886227743, 3.14911376386378, 7.16204977499426, -1.76562842608825, 
    -0.294107989445289, 1.02207973297449, 3.34556285025186, 7.47104260022568, 
    -3.94546864765893,
  -4.04224608315841, 1.31997352189033, 5.52360050497333, 6.85472926555524, 
    -3.31889974420225, 1.50561292342143, 0.235168694870404, 1.37934800144936, 
    2.67458124114638, 7.60797483489545, 4.1958607312124, 0.484992474401184, 
    5.03393685379305, 2.92480416801948, -1.36642059569064, 2.38800083741777, 
    9.91225366373315, -2.043119561701, -1.54934416194132, 0.520072371418194, 
    2.52927862354997, 7.12366364116979, 1.71592897101686, -3.5786246306722, 
    1.2874006787718, 8.03251922927154, 0.864130924754047, -1.55182566327888, 
    2.64529249737317, 9.12713880723929, -2.37558544562831, 0.64534115865032, 
    -0.824786206016828, 0.389319454773394, 7.93719329504727, 8.65610473565488,
  -2.49270138428835, 0.789761515126627, 2.96836138461745, 7.33675467487286, 
    -1.96916629420597, 2.32325160747042, 2.61178841086834, 4.46939828911628, 
    4.86596939362327, -3.54506059899749, 1.28133700813957, 0.556627781029975, 
    5.52864262196303, 5.91609533488423, -3.72436718362055, 3.86948989049084, 
    8.05662453854285, 4.12194514671565, -0.234799950275372, 
    -1.31591943933346, 0.645824223100025, 2.26210061296662, 7.90669544218349, 
    -1.79218695911615, -2.16575866827677, 1.16651895137488, 2.28714443450033, 
    6.2885731277944, 9.08615765542593, 0.0465837237698161, 2.91540763554983, 
    2.6453045238275, -0.40660635178388, 2.64077094395159, 6.87598173632225, 
    1.95949718554174,
  -0.752141351498403, 5.56824212355282, 6.02284150933635, 0.968623339356501, 
    5.33858786875066, 9.15124170618562, 0.432073246128451, 2.84550944514443, 
    3.28367564049819, -2.11920711789146, 1.42132205437878, 2.30985137366265, 
    5.04514121812153, 4.82619425263025, -2.92490874843156, 1.1183444415103, 
    1.44055110110175, 9.28365877095466, 0.212435501237411, -3.25654629300081, 
    1.11620398205454, 8.60976848407846, -2.64576587511484, 2.1249569902447, 
    2.01387217116997, 5.58119860451049, 9.31817065183805, -3.7459122590009, 
    0.110721754842087, 6.38889428251991, 1.72637018893036, -1.04368109537559, 
    -0.538883269153608, 8.10289917359566, 0.340375205799007, 
    -0.285407052239066,
  2.47977674238217, 4.87825061701237, 6.56006465025813, 0.0966424575976994, 
    -2.58051883245633, 1.8288447596523, 8.66925768506919, 3.57654155485097, 
    0.602776727747491, 5.35692873375555, 3.52328624786701, -4.80451348091934, 
    3.13449170849867, 2.53125975651328, 2.53161482100385, 9.12971008289596, 
    6.74308793203026, 0.134707949664077, 4.19444489609949, 
    -0.568124412030171, 0.262184154993072, 1.3182202779121, 3.41637521892476, 
    6.17004494946684, 1.42817375558999, -2.79024083282257, 1.24893744639753, 
    3.13498285296509, 6.66935624184851, -0.869731638746388, 
    -2.10530688094742, 1.38576334551935, 5.59061093058626, 6.02578279963969, 
    -3.69222880122689, 1.91155427773644,
  -1.84813689779855, 1.94666062554728, 6.77798603538294, 7.09645207959146, 
    0.708224341194498, 5.56149978441183, 5.28125775524052, 1.41792932185659, 
    4.32878518365578, 4.15201557845128, -3.33440671401497, 0.969072076722495, 
    -0.0996936132464454, 7.18723411419787, 1.06848619610554, 
    -4.13982164602833, 2.66986714156629, 5.81951480703812, 4.82603557121095, 
    6.22025785412998, 1.34105107664225, -1.14653347850931, 4.01420732431331, 
    11.5183619086976, 3.48864174057562, -0.670941600667606, 
    -0.391596197075302, 0.0723658630564286, 3.28076114950569, 
    8.86916011555965, -1.79047406260071, 3.31016380536686, 3.53240460180935, 
    3.50900991677714, 5.66577507523741, 5.41203439926581,
  -0.524377868647277, -3.34291583124293, 0.502878542243127, 1.3712988834703, 
    7.74468236617534, -0.655872048328362, -4.1658758326476, 1.47711671023155, 
    1.80124243127883, 4.01337577101323, 9.59832257677937, 2.91940516657809, 
    0.295728439347305, 3.12525925623291, 2.049040249601, 4.25021713202094, 
    6.25371372139671, -3.50958176756539, -0.116965579437797, 
    1.66455634324162, 8.11061922486974, 5.54498281054937, -1.56501273457571, 
    -1.56545477006462, 0.365458950801481, 1.31956160948362, 7.98735532804345, 
    0.639433495106178, -1.25683105861563, 2.40515933567131, 8.67709194226893, 
    -0.125010486121683, 4.43991699864863, 3.20347094498722, 3.36459495190765, 
    6.85308954879265,
  3.48593559928638, 4.48281734170299, 7.03629848969532, 3.72763794358166, 
    4.15842241438361, 2.91296850351274, 1.15447871085242, 5.25720435746375, 
    7.82704686251189, -4.09500625512974, 0.889503657447114, 
    -0.349846610521475, 3.79269579062151, 7.39556599390865, 1.96144405606125, 
    4.07625120159735, 4.7775954822299, -3.5216335612207, 2.32834845527134, 
    3.79150034092351, 9.66949154552255, 3.68478160374846, -0.430092353175876, 
    3.09962082321962, -0.949485490685318, 1.6784174701951, 4.78933437084655, 
    8.83860522870468, -3.95815415328411, -1.78280759186232, 
    -1.04615120070704, 8.38696525827646, 1.72071242806096, 
    -0.451993296236628, 3.7514143958126, 11.0434941849908,
  0.689823712142848, 10.058542524097, -1.03343217249811, -1.75728593533096, 
    2.08287310673435, -1.11187020140876, 0.442847684707186, 5.72490460733431, 
    8.63905759775686, -1.42846179951308, -1.2326132734939, 2.76653702485592, 
    7.55831035389381, -2.15907212200714, -1.67749430702687, 
    0.974265431994762, 1.73163987844486, 8.18051005942873, 4.7734768165318, 
    0.276733993784762, 6.31585923019215, 5.17781943126226, -2.20998261180171, 
    5.95803624644711, 4.34954442436883, -0.714922925460326, 0.7030828532492, 
    5.60617024061954, 5.76318231648845, 0.877019508716019, 6.08443050282576, 
    11.2656354516051, 2.33368690653771, 2.3094329983717, 0.423908585650642, 
    -1.67115936835526,
  -1.4900475626872, 0.94452143643103, 1.43258094908841, 10.3056306254131, 
    0.578840503431339, 0.22534650613528, 3.53786212360072, 5.43456354332429, 
    5.04872002963898, 3.92194993291902, -0.907842555756231, 
    -1.55550545110632, 1.72365807244738, 4.26580852521909, 5.30575764270437, 
    2.65088875867586, -2.41635294164352, 1.76076410194463, 3.33285991410876, 
    6.10507879432576, 3.90208809724263, -4.26244107244283, 
    -0.360986591592229, 0.00259824706612033, 6.5712519466725, 
    5.66501831081863, -3.53423535294397, 0.432929793565163, 
    -0.489043973487298, 0.887917116526753, 7.46738770946523, 
    -0.208614008630235, -2.06780882607073, 1.73435355868921, 
    4.24912843713951, 7.53948305440025,
  2.53859945536928, 4.11122265137778, 7.44957410577832, 0.317303489874877, 
    -4.37275513108214, 1.70817658815572, 6.52644188077689, 5.01810014069099, 
    -3.30335275519662, 0.186420973449039, 2.49540228141567, 8.97008032331505, 
    1.95565730329129, -1.86877983098164, -0.449692608328006, 
    0.857391575738328, 3.33739106158513, 8.63874840961702, -2.0622467515353, 
    2.32277401288079, 2.87576206663542, 7.22137242319127, -2.45803046500183, 
    -1.69155661707971, 0.518378449150324, 5.12984951531342, 7.18734398280023, 
    -2.84108910986035, 3.55787432476856, 4.6299066824588, 6.55032019509299, 
    1.79103881879945, 1.71724859068376, 4.88282660906713, 3.03887551264151, 
    -2.86351524298202,
  -2.42052155014384, 1.35244493960248, 3.20077637322545, 8.56789474788742, 
    -1.75398369448407, 1.8154358638905, 0.496748715482468, 2.98109630564428, 
    11.106820190981, 2.97107671926812, -0.267607774913622, 2.34632441982836, 
    -0.645625537872817, 1.92681565132807, 8.77092726685998, 1.5693415143445, 
    -3.04448416593881, 1.29264142210048, 0.873972503425352, 2.3254642149338, 
    7.77717363728506, 0.165613830596245, -4.47275446575812, 
    0.857824249648267, 4.07436987482885, 7.73854253717204, -1.70848452180399, 
    2.51853513164344, 2.4800487694897, 4.06877112333526, 5.6729309159718, 
    -2.72406233914366, -0.0353743287732016, 1.01628678319675, 
    7.77786621064813, -0.739906894798671,
  7.24651723197936, -1.72830127617652, 1.22805133560575, 1.69435626262026, 
    4.80035937388655, 4.93492650543739, -3.51186015815377, 3.05128569192842, 
    2.79067293459698, 3.6475024115015, 6.77702573482159, -2.67756061538971, 
    1.1476837315817, 0.920682657335135, 5.86070324257074, 6.96726483438179, 
    0.449433785017212, 6.19415097553914, 8.76576132680225, 5.47396614642251, 
    5.97500067810803, 0.677513984813601, -1.4419615778276, 2.15010115407688, 
    1.09202289895494, 2.15892912404122, 7.91766590012403, 1.63087065748534, 
    -2.26035691133879, 2.78952159228704, 11.1092799045974, 
    -0.490979757962106, 1.01516618128983, 1.07981839450274, 1.02120894372038, 
    2.96297118380187,
  4.47218756101574, 4.78554501508566, 5.8784128356477, 3.48482673903245, 
    -1.81266373260344, 2.74921545434185, 7.16227157789504, 6.40110949496209, 
    -0.626585236939682, -1.7459426744329, -0.473321030572926, 
    2.06945055218453, 7.28604027244408, -1.10704180265541, -2.44499187180546, 
    1.15789829482928, 5.23979993303474, 8.02502253481101, -4.28383982181222, 
    0.931909950547797, 1.04121327997748, 3.15708054345589, 6.61449880559227, 
    2.37875928438249, -3.3655949409635, 2.87698805237909, 6.23873653015202, 
    5.44332570835069, 3.30034574155494, -0.68421250207197, 
    -0.784609717575203, 2.41623548510656, 7.38101948072696, 
    -0.92466011264964, -4.84792167781155, 1.72100846597025,
  2.26182560504858, 7.83309935317287, 4.72125669387746, 0.0625679294452861, 
    4.75403687045292, 5.65295977881083, -3.83600794954466, 1.46093293384743, 
    1.38328264840089, 5.74446104739426, 4.84215823083191, -3.21928464918802, 
    3.45297761886757, 5.39754608652546, 5.79699546855415, 2.02512565712746, 
    -2.12306526687085, 4.0638325225824, 5.23336879892125, 4.17263692258028, 
    4.94440500464402, -4.34199435917766, 1.15225399184431, 0.777956091143408, 
    3.18176376988717, 8.8669620377614, -2.03765027469793, -1.65223208919543, 
    3.06160836650049, 3.97026230742033, 4.62693341259365, 6.77660787268248, 
    2.4410631572653, -1.30554601294177, -1.66687952956001, 2.08863343432387,
  3.86439463325794, 6.61435571494408, -3.26341803690654, 0.251197485565119, 
    0.685304626850468, 3.33534068152005, 6.57265688407985, -1.10616236454502, 
    -2.00757269507944, 0.614270781387661, 6.63093583902045, 6.26416943241558, 
    -4.19058241073456, 3.113016214871, 4.15149382238019, 3.16468945141849, 
    4.37197793590223, 4.86601303224507, -1.76140960116072, -1.38276395086898, 
    1.30409285295736, 5.73391247679934, 4.10764115864155, -3.29339973150698, 
    -0.686044999361898, 0.707220153904916, 8.61504194023973, 
    -0.408496127262597, -1.92474863638962, 0.28365818450584, 
    3.47842713749199, 9.3825045064875, -1.45009097182657, 0.570188427713005, 
    0.506484568809426, 1.61773921295324,
  1.53197829609579, 4.68800917765765, 8.24338313020245, -0.29591308481881, 
    3.06098726260026, 7.22834185182402, 0.926914717678421, -1.96378302687553, 
    2.76670252177132, 10.1975946959142, 3.53296519214158, 0.105920921991844, 
    0.479162457998179, -0.893669574607147, 1.75548588743957, 4.7852663284129, 
    5.82793657476217, 2.12400853224773, -2.151216529876, -0.606365409193551, 
    1.26089800924003, 6.08407677650491, 5.90547035948137, -1.96197682382066, 
    -1.72778984507365, 0.19617607276686, 2.69932562713995, 7.59932309573472, 
    1.46718795137273, -3.23818769473366, -0.775321793406581, 
    1.01367254443217, 4.44954976734061, 6.70605948793459, 2.06549163789108, 
    -2.77451357157462,
  3.37476697107564, 6.46596936304515, 4.32961792917742, 6.37924998475977, 
    3.17922988079746, -3.26431492793734, 3.40527435451246, 5.67216906118077, 
    3.26430400530788, 4.61013399677506, 3.3651600970444, -3.54773861712752, 
    2.09636397299422, 2.96710852553329, 6.61607656205651, -0.216854901862386, 
    -3.94551567436983, 1.65367500821388, 2.43560782098163, 5.01309221738135, 
    10.7945610026853, 3.75187561050224, -0.189708622719926, 3.30326635924778, 
    0.00392400493395018, 1.59366935955843, 6.85321871026909, 
    7.07520530399317, -1.77312391496832, 4.76403159889007, 3.891523780605, 
    0.548652411729354, 2.5558202520626, 8.60534959628599, -2.49240463306313, 
    -1.32672741855929,
  -1.27057341445356, -0.0899605201188312, 9.09668185995477, 1.08412510777114, 
    3.68309671929914, 2.72694458070582, 3.88226492351764, 9.41187687692023, 
    4.31017624047294, 1.89919283618944, 4.86546285601198, -1.10031296236192, 
    -0.733272608061814, 0.760045570984747, 2.48461021222884, 
    6.78174959960527, 2.87102561933313, -3.95698894559954, 2.34786651677196, 
    8.51843332007491, 4.95331529975923, 2.48330794765874, 4.13410775430611, 
    0.316800328554027, -2.13989320054914, 0.728193019940212, 
    2.62129635061195, 9.05272006278093, 1.19104823847572, -4.14141781457797, 
    0.744374696288565, 9.11095571688967, 4.91481107649928, 0.127707815923015, 
    5.25328294003549, 0.717102887905685,
  -2.67718667338911, 3.4429463101797, 4.79360020293443, 4.08084301099322, 
    5.43374479690869, -0.156308246925747, -2.79290849827914, 
    1.51876809640239, 4.42560901249401, 6.17921102615069, 2.05676484742294, 
    -2.9490513523328, 0.294933248111144, 1.93770004163148, 6.49558485287181, 
    3.28643302530599, -2.95492608382498, -0.136818923948566, 
    1.48897449892299, 9.27407582178159, 7.07447509810255, -5.72796954840168, 
    0.177606143076201, 4.49331940055627, 3.09530903054584, 
    -0.877776500214818, 2.41737016623029, 10.4575676192493, 
    0.839479660642439, -4.32389898197716, 0.028005525072015, 
    2.97575682243639, 6.034647145569, 4.79304945486811, 4.86919558312268, 
    1.90831923707659,
  5.18385411589375, 8.62010507941047, 2.05466003874167, 3.72063300617864, 
    2.58846213807607, -3.40128318361371, 1.41920036874004, 3.12853959807809, 
    7.41056084531861, 4.89763065551675, -4.35013724270715, 
    -0.761800867818527, 0.551172796220509, 7.25276275313664, 
    5.77152794510111, -2.17997653633194, 0.0390330572010313, 
    -1.15607893762528, 1.41056947941038, 6.82997471481855, 5.4149142136508, 
    0.287320229846494, -1.00688460322128, 0.1317165051202, 2.50300852172843, 
    9.70496835307669, -1.39730844811696, -0.0959305717735868, 
    0.732469558631008, 3.3757719744489, 9.08481676243094, 1.89739411790217, 
    3.73318589446964, 7.76228577387242, 0.547272794108628, 0.685510674376402,
  -2.76099465370116, -0.661629543455777, 3.21908721216398, 10.5188141295456, 
    6.88873487209151, 1.48533010090692, -0.0256195969741317, 
    -0.394467791679341, 1.49924871569451, 6.8892571694477, 7.89077798554302, 
    3.9360986280949, 1.93962958955514, -3.10931367519839, 1.58495514956075, 
    5.72773286851689, 5.95921020993136, -2.38189441474441, 3.1909537358863, 
    5.87247087930259, 6.39080205003372, -0.459377810933981, 
    0.0457409904565522, 5.00568504803785, 9.41081858957966, 
    -0.455178941627685, 1.44419593664269, -0.670332835523283, 
    2.13692129581955, 3.73195257249934, 8.62306283102728, -2.13552582819692, 
    -0.566013701118032, 1.68790594384695, 7.66085800951344, 2.59905802604965,
  1.56893557606515, 7.47611006346542, 4.15927982708063, -3.92429593616258, 
    2.55015861686891, 2.90240962147535, 4.90323366934525, 4.16640940138023, 
    -2.78788008980972, 3.07212281603955, 4.1788412594657, 4.40872265687674, 
    4.49351106211591, -2.27642525579777, 2.53931663186951, 4.16569084165247, 
    6.50712416493003, 4.55987155125286, -2.51518778139724, 
    0.0237943254846726, 3.2032668121633, 8.71596447817442, 
    -0.105459846908143, -0.722780534354798, -0.290225966928032, 
    1.67880447583074, 5.5143175161396, 3.97718452562027, -3.79735052361777, 
    0.898970830149968, 1.47432239087819, 4.45194148979528, 6.30381544529114, 
    -0.945890926964324, -2.96588613284269, 0.743537338440408,
  9.87934217052771, 0.7183758555531, 0.992182830000576, 1.86095837397079, 
    0.814799492577451, 2.86956183966719, 7.47959197815032, -3.14465687407211, 
    -2.96546750822074, 0.106770015115657, 4.28258007312231, 8.10769597095522, 
    1.30457828611717, 3.16484302459775, 4.27908494133136, 4.19485357121356, 
    3.11642160711398, -3.34249462042882, 2.20810536034663, 1.56666662554398, 
    5.9775521365388, 9.02168033397804, -2.10767310349947, 1.08331877919065, 
    0.499619970829917, 0.718846209489285, 2.05563608435225, 7.08845513874048, 
    4.48390116890684, -0.492700844952263, 4.76120637236146, 7.6526544330693, 
    -4.07731033992194, 2.63293702827611, 1.16912685708903, 4.12772919724345,
  -2.64226027263152, 3.64628304610812, 5.97329022406663, 3.44084759429071, 
    3.63844126226117, 4.27866850477186, -1.3310957904189, -1.09470782663114, 
    1.31451625992756, 7.70401067310136, 4.1544975895329, -1.46682749062785, 
    -0.806960218837351, 1.41530691675342, 4.0737034600106, 8.15260124586875, 
    -3.61808284377582, 1.53898274856651, 1.61482608284389, 3.22451357183458, 
    6.43106332675828, 3.47395372608561, -3.9279951211289, 1.86051345295712, 
    0.289463929418892, 1.10146469311641, 5.15675656914813, 9.29761863402916, 
    -1.02012161366028, -2.30946550282802, 0.942830274908246, 
    6.61511309416942, 4.14611408449551, 1.12486252550259, 5.52220059445097, 
    8.42261073529104,
  5.89915788377771, 7.94922119590546, 0.803726608525451, 5.17627618719371, 
    4.46453058277661, -0.236884535777902, 3.83192983219609, 6.39583617205937, 
    -3.21441380975513, 2.71108774502039, 6.39703186211253, 10.1104383270678, 
    -0.807015702716893, -1.87337793648612, 2.19680823190983, 
    3.28514266998484, 5.62949896618763, 3.85275523559338, -1.61308651053269, 
    2.57048618694871, 8.6504266396899, -0.20549262677349, -1.44311240372845, 
    3.47157447809512, 8.79771001200386, 3.34209170511459, 2.60930585856078, 
    1.24116842834287, -1.77689873449337, 1.49821638213098, 3.10034385264274, 
    6.08151798471565, 2.53829559140397, -4.74384844191426, 2.70209778367126, 
    1.54736365157588,
  0.522315585059741, -1.92302083414017, 1.85587410245599, 8.01048170885465, 
    4.28007595014943, -2.67886150308004, -0.773563608230324, 
    0.624455769903782, 4.38042200572445, 6.96785195798508, -2.68493560185367, 
    3.72899419359447, 2.42104845058247, 3.79228725677201, 8.12347390411076, 
    -0.781382536376354, -0.747440229300363, 0.791566290048556, 
    1.92678440310009, 4.28181485957306, 5.73243076364019, -3.44708329975146, 
    -1.29483027717276, 0.0215801713711703, 2.1322628403575, 6.40471994287332, 
    4.27323578762693, -2.72680723141268, 1.92271004706652, 6.81552689010053, 
    7.62511112817028, 0.00521936490499986, 4.51812769493545, 
    7.02649778535741, 3.76651472168262, 3.21512427493366,
  8.09213100273708, -2.29346461919057, -0.121977757059657, 0.590692065396532, 
    3.76750575172315, 7.8454221843822, -2.16560279213654, 2.47996131755599, 
    2.13271815416843, 4.67540036829716, 7.91740539466015, -3.59861580421488, 
    1.7844997793798, 1.43075421883654, 4.4771867167935, 6.35096635063727, 
    -3.81938941168943, 2.58421798081215, 2.58793313323919, 2.74866424338452, 
    4.39557675803262, 5.1724964134913, -2.91279813932416, 1.68424178343443, 
    2.61232325316011, 5.32872283487717, 6.92629184052214, -2.14087162192571, 
    -0.682788232618399, 2.3201558698817, 11.6487563164449, 1.26054230589623, 
    1.58759288928132, 2.09082268186844, 0.716313122174242, 3.18962513233167,
  2.28827343719095, 6.08903594934693, 2.54067976428572, -4.65459407576042, 
    1.54664276153042, 2.28765704548681, 6.14779319485323, 7.75579745938727, 
    -2.87307004372796, -0.72710299441939, 4.1193477253803, 8.20331865038579, 
    2.759964050876, 4.85466682282937, 6.54340147247814, 2.13910605669104, 
    5.59257095260399, 6.23873623392898, 2.41392252214448, 3.63516829808056, 
    -0.255722690567753, 0.423343315035612, 0.477126073633751, 
    9.02964915990739, 4.52280872269689, -1.25424730361577, 8.2461693678396, 
    3.42344621087069, -1.98157597779091, 1.32481054154227, 8.09395148573568, 
    5.80241142673305, -0.64405590162396, 4.24828121570587, 1.93449946610028, 
    -0.31953166679942,
  2.17834820007832, 3.55076866548607, 3.83821712996722, 6.94021484570783, 
    3.59777811400833, -3.60997502171737, 2.99776717191182, 3.70018565605069, 
    1.58103709842413, 2.87997123131874, 6.96272613752415, -0.738566922957859, 
    -1.58255149786938, 3.28131288868897, 8.25440500185661, 1.9709571863382, 
    3.97866654563032, 4.84655692323137, -3.24176792389488, 2.07230504608243, 
    3.76595564151078, 7.50333805601295, 0.667588019441917, -4.24216140821797, 
    -0.0371195517621281, 1.22686832902322, 8.37001206271198, 
    0.0567787084334204, -3.24650665086416, -0.63374783760071, 
    2.24376650014631, 9.92336097131114, 4.00429025411327, 0.123835909971134, 
    0.403865137447718, -1.44432520085389,
  -4.31752612500864, 3.19331974514254, 3.20814445296426, 3.91703807723569, 
    4.60575770218534, 5.32242885583027, 3.57217210757462, -3.35518262209846, 
    -0.651941370182177, 2.26097373843742, 6.8564355141557, 5.30442221636417, 
    3.94473216483128, 0.931213059424899, -2.60002746028728, 1.81842097685392, 
    5.36099628237105, 8.47979596796193, -0.332879828988861, 3.61715502166896, 
    5.96361210334848, 7.53369582421757, -1.48473069913493, 
    0.0595831365972379, 6.87718622036091, 1.84443892203621, 
    -2.96322118784088, -0.73249350129507, 7.26286217134514, 3.79839381360435, 
    -0.357413759927651, 5.92229413230116, 6.93206791574784, 
    -1.60617548366136, 4.49729173842223, 7.05024724077621,
  3.29300647466333, 6.74724099936992, 4.22915367956151, 3.74739803224085, 
    0.735006348301945, -2.51444025216327, 2.31083944302239, 4.14189773043736, 
    6.49776761958207, 0.246151913422293, -2.54121807477828, 2.6934690894664, 
    8.80076452874531, 1.45280748077802, 3.48977144520779, 5.49173271476946, 
    -2.29259000221181, 1.17721725756335, 3.55281536170766, 9.1466114312778, 
    -1.37984481184601, -1.01520347638888, -0.82253488850424, 
    2.33553344629366, 8.08086571312826, 0.756192276095249, -1.60228972772821, 
    1.32525982845063, 3.26522599094182, 8.57942818165384, 1.43154940634585, 
    2.08892962517246, 4.48394780224588, 6.53177783085803, 1.27169224182952, 
    -2.43452638854418,
  3.92871693712765, 5.47456843652987, -0.752563934281833, -2.03323222414967, 
    2.76269932216701, 7.53117538704382, 4.57047342122263, 3.61227526942731, 
    0.352373081246754, -3.27130557006675, 0.992299823011761, 
    0.150364830272707, 5.70978158747512, 8.93174856988486, -2.32250193323999, 
    4.40995261273199, 5.06171626852728, 0.399624726439384, 2.32747479371113, 
    3.98325824244355, 5.49040466394361, 2.51951908094555, -3.41372255137964, 
    1.98964781343051, 2.03089729376402, 6.54113203473186, 7.44813778757241, 
    -1.9459861079714, 4.37022256712348, 8.33830224701322, 4.6332262997111, 
    3.81614195589956, 1.05390879324719, -2.1064821628806, 3.32127594959235, 
    4.68601710884667,
  8.68969713989854, 1.068642958529, -1.78883506526439, -1.08186253064522, 
    1.94096922487921, 5.51562558319941, 6.39098101715746, -0.371811023192643, 
    0.522890824758801, 2.81313027713659, 8.17388303595873, -1.73771576781491, 
    0.176055971790006, 1.24974264111783, 8.76728313412411, -2.75383365249192, 
    0.352073915871039, -1.13863997537851, 6.89699560422375, 4.72246873711759, 
    -4.33540121082492, 4.4754395118979, 0.844433839235523, 1.97764207236246, 
    5.35183825438241, 8.05332613748095, 0.833138027923911, 0.882857897746816, 
    5.73777440156894, 3.15598135776821, -2.31366216952918, 2.02566057022011, 
    7.25773989614847, -0.138257472779523, -1.46289093413575, 2.0755077214998,
  -0.861388922109034, 0.191657559643713, 4.7902754574724, 9.39888198658122, 
    1.11799656539173, 4.17368862510348, 4.40241682648905, -0.294153971162235, 
    3.39138169464306, 8.43658519514631, -0.430014799266707, 
    -4.96281413629219, 0.994679199915837, 5.81703316120989, 5.85798997366299, 
    -2.27511531412315, 3.93730863727341, 4.26522855468193, 4.99331846940322, 
    7.02706063634297, -3.13396434878211, 1.26276928409428, 3.04031376540415, 
    4.40416359516762, 5.2973506036959, 3.93909916759437, -2.70233009825617, 
    1.16679534888427, 3.38434097069008, 9.51245887949363, -2.0036083845864, 
    0.301654380110869, 0.773378074802542, 1.98050973180173, 3.93536916296728, 
    7.50700588737723,
  6.57290124722143, -4.8077438962551, -2.81784553882764, -0.481666994196568, 
    5.650908648314, 6.09634971957827, -0.99126485372329, -1.45623592593955, 
    3.23314903620341, 5.31285921425918, 4.97059174368961, 7.44794275693797, 
    1.42084476718088, -0.218339240343154, 5.52966960900176, 9.02333596513108, 
    0.478935536629189, 4.37251214857677, 1.48636902235482, -2.03603513692483, 
    1.55043303271929, 7.07606418674829, 6.24380807570349, -1.28315109953923, 
    -1.18762268455801, 1.31067220833273, 7.47323194610225, 7.37622703441805, 
    1.31109068914284, 4.79714590325681, 3.42221728433681, -2.79521017277585, 
    3.85795322575252, 2.142629648621, 1.48313499522898, 3.48712708826604,
  -3.59626787270387, 0.803303933093915, 2.19468391328148, 6.12066081855812, 
    4.81868665191465, -1.93358734264756, -1.52959249484108, 1.32443203824258, 
    4.75100496845952, 6.46110745092029, -2.64180353722724, 1.72636971958653, 
    1.99270309616888, 4.7195901385875, 7.41949548457118, -3.14900933786292, 
    1.48749778189537, 3.1709968322043, 5.51544245718, 5.31640848336309, 
    0.334679042893216, -2.77733062239384, 2.69240930203462, 6.43216626759676, 
    8.26883620865829, 4.94348757086502, 1.42879081022378, 6.30691992085573, 
    6.03648856417573, -1.8155965922727, 3.23250564732916, 1.16306905384525, 
    1.09554766604809, 2.65928624534491, 6.03501362785599, 3.00447806472555,
  3.00289956267776, 8.4063825743462, -0.359167064502519, -2.48933509217103, 
    0.450660599720923, 4.0545765303932, 8.83282425139756, -3.02130621942384, 
    0.85376918247293, 1.40911963488995, 3.06617801885733, 6.97689807449966, 
    3.07762870095129, -2.33746351380795, 5.45098597177943, 4.13156527430711, 
    2.22157460535277, 5.10477931451172, 3.87649023393935, -3.03873101669233, 
    2.19360632613391, 3.25086521572494, 6.70771939590326, 1.97851241986498, 
    -2.24963041860214, 3.2754758193144, 8.24356889687836, 3.36462658074559, 
    -0.41686221355205, -2.07232321965643, 1.04984919949182, 3.32840231858392, 
    7.32053695692788, -0.935077821421963, -2.15136866499748, 0.38322986432369,
  -0.726440154383914, -2.12819148286185, 1.48580766073948, 4.72721546070268, 
    6.56797349948239, -2.40326443516051, 1.95067731492175, 3.34503713181831, 
    8.66784345790791, -1.94610698674944, -1.77609727680853, 
    -0.143466233531705, 5.58651586842206, 8.5664185266406, -3.70720348939488, 
    3.95900415066279, 3.29820033137176, 1.9823500264566, 3.68299209159313, 
    6.22512143825825, 5.53184467991363, -0.11063489511965, -1.96760014112834, 
    1.01077797580353, 5.6592883609829, 7.00514983260791, -1.70819625625365, 
    3.97725588656187, 3.69848624349159, 3.74383233875581, 5.43888519712787, 
    -0.554815978688628, -2.35910548021068, 1.67765517935773, 5.8091345966538, 
    5.56249091987419,
  -0.918607280913673, 2.49845633190998, 8.91374464547051, 1.06560150380297, 
    -2.99365024352531, 0.0234139545402958, 2.37648199877069, 
    11.2501467706723, -1.9925192343634, 2.24241346598902, 0.607003516071526, 
    1.08354615812777, 7.51038201553182, 11.131077369406, -1.09848246824342, 
    4.24576925263603, 5.84417770743504, 2.31508463875476, 5.03619202255902, 
    4.23755740605306, 0.263181153732889, 4.03030092551348, 8.39462113866175, 
    0.251307810678235, -1.75484602443998, 0.11726268040341, 1.38609654823569, 
    5.09146663245409, 6.79884884111223, -2.75175739268126, 3.63647590842996, 
    3.57914673348871, 3.26490847709581, 5.21198484621434, 5.22679134872693, 
    -0.828897110679106,
  0.133497451451155, 0.786108245054174, 12.0263292434396, 1.95628401890959, 
    -2.32655607075656, 4.0982201923792, 3.26006684003878, 2.18131607722343, 
    2.60437611710927, 4.01160427989505, 6.4206579816685, 2.19963474516784, 
    -4.1780139675616, 1.61840760418554, 2.53984814386497, 8.64728985343522, 
    1.76583056438035, 1.5976826236, 6.37681137491532, 4.69520057533676, 
    -0.752678854191358, 5.90527725544062, 9.97645234199352, 1.99525116487839, 
    3.14899923224094, 4.24334148112009, 5.47821277831188, 3.39537351881231, 
    -0.630963719364967, 3.52946559573352, 8.84363876633145, -1.4943304180061, 
    -2.36289112441325, 0.736407402496163, 7.61837507764406, -0.951552712249328,
  4.91205105183666, -2.64450252814127, 0.579900551457288, 5.35076473753151, 
    9.36012476688795, -1.06447286064622, 0.19954074966477, -1.37441775834984, 
    1.36974192851283, 4.48193777975105, 6.58264587202677, 3.49440429001375, 
    -1.51135552027883, -0.66584773245624, 1.10545288746217, 3.82292084250049, 
    6.52249443352423, -2.26322440542762, 1.48439767292877, 2.36268907784695, 
    4.50443311051364, 5.25067099705526, 0.269465428840825, -2.88624175860418, 
    1.05932376348316, 3.20567545341167, 6.65048842820255, -1.52125693801781, 
    -2.0079896038049, 2.558223227057, 3.79035825628665, 7.94666106879455, 
    -0.516762830739507, -2.70875312482212, 1.02698001784085, 7.88351358162914,
  2.16075375105734, 7.23294249687059, -0.871991909793731, -2.57539819410347, 
    1.56876638502403, 5.22624870792902, 8.23791847733419, -0.426911763264416, 
    0.948601281586639, 5.60027864956088, 8.02872752997948, 1.49039559653162, 
    5.18965339502696, 8.13932473441315, 1.94672015582197, 1.71045850114057, 
    0.388064493810101, -0.396731223680916, 1.743290609608, 5.91020437688169, 
    3.92640636886583, -3.70161780671781, 1.30868446911307, 1.68381292867352, 
    6.63237969158423, 6.27155770808673, 1.30065267242257, 6.09100761900397, 
    9.89513165098686, -1.17604750552689, -0.0891542619672827, 
    0.178259750311316, 1.8139927074709, 6.15758480051861, 0.0174767964817866, 
    0.266043014901429,
  7.97339008159125, -0.32997430203204, -4.70304066946885, 1.90506491982157, 
    1.16129368087504, 7.56443870898197, 6.68265504087539, -0.191545212333295, 
    6.76432139722299, 1.69949046958577, -0.796177987508618, 
    0.787280043957756, 8.87385490146518, 6.50779204776245, 0.589451226512242, 
    4.28756501461931, -0.788226379855724, -0.428112999191179, 
    1.54248656337698, 7.91208162399439, 3.05378154979103, -3.86852642886954, 
    0.176284532413328, 1.27329505815794, 10.0336888906058, -2.19016645971426, 
    0.356114881469469, 1.20095857297798, 1.42547166234432, 3.17721185605633, 
    8.42222062752301, 3.59144143892736, -2.22211382036684, 2.00393200706232, 
    0.794824949426191, 2.48342701228622,
  2.41101025883435, 3.29240856730906, 6.3075441784429, 2.82538679465223, 
    -1.78167797185148, 3.51079085800481, 7.38645131571688, 3.50717771716645, 
    -0.907617428037532, -2.50381817232074, 2.07117655823551, 
    5.80618598930429, 5.18681081900043, 3.03529377180374, -1.04915869153475, 
    4.75669104826712, 5.88545670817842, 5.95077332876504, 6.99366384257606, 
    -1.21465148782386, 1.97623565691144, 2.67248559007464, 1.95913369362178, 
    4.60730280432163, 9.1472236461453, -2.99750133381597, 0.088906963528693, 
    1.61062983394448, 4.67964049361673, 5.39194515102325, -1.21367298786896, 
    0.256538921937859, 1.89966494032267, 8.97965172863926, -0.1650802476451, 
    2.66197789032962,
  4.35583955513906, 5.9247422876377, 1.75241252449681, -0.838577021957128, 
    2.93809152574877, 8.67935594530984, -2.42638411079195, 3.11456909879802, 
    3.3723911710443, 2.34140346851114, 3.67915459387365, 6.20353309620735, 
    -0.156477599477277, -2.55745834034136, 1.78496769593022, 
    4.77939968591536, 7.04368082825824, -2.43514082878219, 
    -0.386978089408945, 2.44047404154507, 11.0938602496112, 2.87048677177441, 
    -0.145400631962031, -0.437462733318009, -3.63901620264839, 
    -0.36617950949398, 5.88646601689317, 6.4604093652708, -3.21910932804086, 
    -4.70783237679894, 0.227287867134892, 3.12739799973861, 10.3547631240296, 
    4.84644937487446, -1.66129321909131, 3.00038058122996,
  -3.38391601149538, 3.61315720558881, 6.57476386452787, 5.26069150845116, 
    5.43652365391972, 2.83352593181143, -1.0284922446629, 
    -0.0912826701979896, 1.13681503451363, 4.65342720406047, 
    8.05360881408009, -4.90564446447111, 3.16957118526655, 1.29402079604174, 
    6.44471903074372, 9.0062318582825, 1.15439576371854, 4.10652374872389, 
    1.90724189271313, 0.257854297531515, 4.61428114138645, 12.0115881701583, 
    0.407240872058105, -1.34112698439831, 0.278196586185754, 
    1.27902374169388, 6.1455722882776, 1.74913025236176, -1.98456891109975, 
    1.08753490019258, 10.0565745038957, -0.0563456827410187, 
    -4.4324801364039, 0.237651854611542, 6.19389532123339, 3.7768709561153,
  4.65782341089637, -0.765974832511061, 4.23988243647425, 8.91520004550563, 
    -0.83219648884996, -0.944016760377225, 0.193057745627654, 
    -0.311673037104183, 1.00314878136382, 7.67051497077203, 3.8944148618574, 
    -5.71590602493609, 1.04398812313176, 2.11088808770022, 9.51310488698386, 
    -0.504051580893186, -2.0829680684101, 0.909013120047398, 
    1.03074209386331, 3.20193299197786, 9.30343780558085, -1.53119222883146, 
    -1.53025788662814, 1.25392009767113, 3.48894830498602, 7.00517142732724, 
    3.42622181644243, -1.66243693302914, 4.54866936066595, 7.78686189516956, 
    4.07008746405994, 1.81739715398014, -2.31355325629604, 0.796018948589148, 
    2.08661560391826, 7.19074909956343,
  1.2773339238768, 4.64851532525208, 4.63629668331204, -1.41678448141115, 
    3.64049296942113, 7.5060470072148, 2.08985383998778, -1.45988599794722, 
    -0.953716790035099, 2.16235740118451, 8.60366054006558, 2.94332170407539, 
    -2.90845257884692, -0.788285719384813, 0.897635318899235, 
    8.2383750433159, -1.15121675976609, 1.43497276104725, 3.68436497219477, 
    8.96011555701151, 3.41421456102967, 1.45996589046398, 2.51294235470828, 
    -0.587673251247803, 2.59167307785608, 7.07111748166495, 2.41605364470427, 
    -5.50080461622692, 1.44241488477375, 1.92233743275666, 5.64173204198628, 
    8.80279447469848, -0.411059622638186, -0.425951899768081, 
    5.23793339890576, 5.24618013620569,
  2.19369677600617, 7.13400313406135, 6.00700871062668, -2.89234410891777, 
    2.72525750928746, 3.1704589671376, 1.04151681933364, 2.69930873083494, 
    5.61600190442741, 2.55000704062369, -3.48525258570621, 1.75456702849243, 
    3.29789678438537, 6.62308374053048, 3.86225150477801, -3.26130996462851, 
    -0.183113329740296, 3.12133746163743, 9.76224410145333, 3.37592835458394, 
    -0.671563250599803, -1.39238402612886, -1.43768188694165, 
    0.796009421717281, 6.33215131473559, 7.34496298961584, 3.18330475051506, 
    -0.415630878389417, -2.7392042405735, -0.298334280242348, 
    6.61585336427601, -0.0707455236777963, -2.80822116254684, 
    -2.46295107053335, 6.97625121428783, 6.44066519394366,
  1.23866150764891, -1.22813379215547, 4.7974398541628, 6.55477186641346, 
    -2.46465255582032, 2.43619487894695, 10.4657755260041, -1.56156839683657, 
    0.298766225464301, 4.76815093549965, 5.6235743535094, -1.76923128677479, 
    4.30908775318724, 5.87243836215056, 4.62254227763863, 4.30815984530967, 
    -1.94164971966332, 0.631705009158508, 2.71191372912654, 11.3465373103481, 
    -4.1341292159311, -0.28230623430859, 0.0723114694859119, 
    4.39177433006691, 4.84518220720336, 1.33197998074604, 4.17212401456904, 
    7.11597074764412, -3.43321371664465, -0.270113420835922, 
    0.139629429052708, 7.13568332861867, 1.61323301893453, 1.15410861648873, 
    2.35274287180254, 7.35674674648942,
  5.54738288630607, -2.7688405439894, 1.90699533107382, 2.44248843089839, 
    5.00849474104828, 4.24140822446328, -2.8873719020418, 0.538628260503427, 
    2.26403401245879, 6.47488030972798, 2.45428220907865, -2.3073065547883, 
    3.0381141939305, 7.08354802060481, 5.48046443239079, -1.6551085452701, 
    -2.41606191865114, 0.979092938582016, 2.91934374105927, 4.97099308306125, 
    4.5837772184436, -2.99563982350131, 4.70800100459639, 3.67674051865121, 
    4.83435294392563, 7.15660518684472, 1.19610541084357, 4.75874239163947, 
    6.18433078809495, -2.55586043147475, 2.9292883864789, 6.38702223147261, 
    3.72550357022581, -2.40754854761366, 2.15731424590972, 4.87212536716216,
  -1.23970121882304, -0.810548625748868, 3.78531903021261, 9.54760465808957, 
    3.95028931298172, 1.96202565968117, 1.02096233197241, -0.8663268830908, 
    1.53679665071249, 6.59553797559543, 6.41490381846051, 1.24630313465196, 
    5.53089401892839, 6.67459620494056, -5.16485206046631, 3.71931319873835, 
    2.37813725244443, 3.19474363230324, 2.60802492124498, 3.92495831408744, 
    6.76250022006711, -1.16925872955921, -0.784024079511473, 
    1.31992029580598, 7.75840457972008, 2.3078646303789, -1.73459337876665, 
    3.4039771714888, 8.86311736469353, -1.97674758911947, -0.523240470136233, 
    0.0878173905059478, 4.03515324793631, 10.2700843387222, -3.4666433926352, 
    0.260216570976237,
  -2.53422130475197, -0.789846071019755, 1.28128261198375, 6.4417033890349, 
    4.01411834395839, -3.78778373917225, -0.824721412339638, 
    -0.45400342194234, 9.1428071261738, -1.85107911746922, -2.04219769163458, 
    -0.312572589578521, 3.5427987034538, 9.15037545558499, -0.87472579455977, 
    -1.20870633216666, 0.87138702507646, 1.0638245145023, 2.34986360153693, 
    7.48859346186791, -0.479987663569326, 0.0739387606207136, 
    2.16955622120881, 8.49905612864961, -2.13944042070712, 3.05195439246316, 
    1.44008110531711, 0.401188116929652, 6.3642682006135, 5.51355670566287, 
    -1.24871407584424, 5.85056127588465, 5.70089835018314, 1.05252196313274, 
    4.07697435578738, 5.41042474889663,
  7.98756856636693, 5.75966350741084, -1.25007688141678, 4.96644700317263, 
    5.33421349301822, -3.41585672500042, 2.59014707362566, 4.17244080911635, 
    6.93278218914151, -3.62910110163479, -1.16919678887468, 
    -0.941231629498977, 7.60868430530906, 7.59629582938885, 0.86553824455695, 
    2.06238478568475, -1.59668454085243, 0.87441837138061, 2.04125563860439, 
    4.48026804303912, 5.90989462076627, -0.339537236252673, 
    -2.10291540429638, 1.91779222697697, 5.10991202691541, 8.65135130188659, 
    2.11370113824835, -2.49828402852759, 5.8670293919717, 5.06875054346649, 
    -1.44518733175253, 2.57416971403725, 8.50502841787148, -1.17712052137226, 
    -0.648569069596826, 1.20205435424692,
  3.03385090927988, 4.70857709053538, 0.521316442825004, -3.74055688941313, 
    2.04960227345453, 5.08069215832987, 6.16485142258659, -0.277134944990623, 
    -3.1362146782611, -0.236013736528335, 9.30432793108934, 1.41048720151655, 
    -2.80674769759801, 3.78376367618954, 7.79594365010312, 2.35773855932749, 
    4.00073510222151, 3.62024361815332, -2.82569798115706, 1.35150119351056, 
    2.56304109353279, 6.41772140323445, 2.00750916947072, -2.82354990000106, 
    1.05547002926522, 2.53093815124593, 7.25033506183653, -1.47289891168146, 
    -1.39495788022271, 1.42153558234896, 8.05580545479491, 5.65945750468204, 
    -1.7669468574196, -0.336789737054445, 5.19663300308292, 6.86088377282749,
  2.53827104995441, 5.23071927958604, 8.87608260375028, -0.926414283960516, 
    0.754841087539675, 2.5394237315003, 4.29386184832431, 6.73855046899966, 
    4.735612204418, -4.86456163871056, 1.08804558797743, 4.67707182384271, 
    9.17845153589906, 4.49997948450318, 0.286747290342608, 
    -0.775973594352738, 1.79519313532475, 9.41167839284412, 5.29195784117311, 
    -3.61747250827646, 4.67747400834225, 7.55856275049474, 2.57707694212501, 
    4.18689677613304, 2.64602971108073, -2.08047489308524, 2.22828246331994, 
    5.00776586536427, 5.05476592179838, -4.03677779966366, 0.698428705098502, 
    1.19753671871408, 4.65290717260782, 6.3815042580086, -0.0710445361697207, 
    -3.49569853548709,
  -0.519560725031043, 2.13151421156626, 6.29377778807178, 6.09699079380416, 
    2.29644130488976, -2.24861304544896, -0.685940113720195, 
    0.594087846733988, 4.37194989275258, 7.73752645520602, -2.74729351918858, 
    -0.392775249841062, 0.847707832039757, 2.30024195386276, 4.1435312582535, 
    6.09286516946503, 1.1576568264991, -2.30768942887023, 2.12484630099398, 
    6.33016201336986, 3.45915678580273, -2.86167099076638, 2.42415534857312, 
    4.68629508759816, 6.3630020534177, -2.40713228905463, 
    -0.0784545454441283, 1.03648851057718, 7.70942593186232, 3.0627332470093, 
    -2.36035817887556, 4.1954173665549, 8.96859564729614, 4.1609013467741, 
    1.44196686860972, -2.87958099397059,
  2.52806631816613, 6.77792786746949, 4.5373690346034, -1.43069135774603, 
    -2.4276843328541, 1.00311181240833, 3.74492336384283, 6.60494348322961, 
    3.54946159911013, -2.16004505445588, -0.890087872057416, 
    0.878572646731583, 3.21642975995685, 6.78250947497912, 1.50757759703581, 
    -3.13967483231654, 0.862592176528326, 3.12321860587841, 7.38976799531825, 
    -2.88491364148593, 0.998442823157569, 1.79245023248859, 7.04873850491954, 
    7.44313636424141, -1.56966839731543, 2.65275614694365, 7.1847216942919, 
    2.79931374375686, -3.58118998704018, 0.548343769473471, 3.29515698070072, 
    10.5104405822028, 1.20763737127733, -0.561494945519099, 1.58465732055915, 
    0.0265715908806423,
  1.1815323536761, 4.12909972846813, 6.2042526045581, -2.2172414169092, 
    3.00116240325285, 3.62381140782755, 6.22755876526241, 1.95677350565367, 
    -3.48387185429912, 2.40295339029011, 2.64416869048428, 3.97100136531971, 
    6.94764965438685, -3.2939186586503, -1.11920639623023, 
    0.0142348612786156, 2.85929712856724, 9.39923309439688, 
    0.665346889709317, -3.13397950233343, 1.83445387083302, 0.37556481681736, 
    1.01695266170143, 8.22608470363325, 2.08165357034234, -3.62127101021334, 
    2.87329580832014, 2.75045793415962, 3.29495556066455, 6.52349457014077, 
    0.744481454162483, -1.63852398162349, 2.38650910950744, 8.11110449551318, 
    -0.459676965547073, -2.05383037781936,
  7.55843139932326, 0.612808551954959, 1.05639895389188, 5.49488614191219, 
    3.92358721025011, -0.3380420320111, 4.08983529007221, 9.16017068363672, 
    -2.11817719205984, 0.366675170794462, 1.51823738825881, 6.91863065322382, 
    8.94324662283232, 2.41168415939037, 4.85535572239291, 2.93786282006615, 
    -3.67345280224357, 3.03045472176906, 7.29727983740656, 7.75314718100599, 
    0.514336322887498, -1.90258835434716, 4.39045558063515, 7.45296168730771, 
    3.66558547322775, 4.94754903724555, 2.02630829312922, -2.18637809116611, 
    3.74228996155346, 3.14777838042951, 2.8634844896909, 6.8523694760232, 
    -0.608408886221098, -4.26878224327015, 1.42476284839576, 5.41624257242449,
  3.18102538484665, 7.30849753681852, -2.2971024577611, 0.00641172829641334, 
    2.05203401675749, 6.03353607372206, 5.13780547073711, -1.54582523930682, 
    -3.36596254026931, 2.42210669788271, 5.33878080004832, 6.27914453458941, 
    -0.593473428337847, 1.28187997260925, -0.0810949013518751, 
    5.95669783752919, 2.89544238190529, -3.15088734458787, -0.92498904177962, 
    7.51256446631554, 6.55762456927628, -0.153515147729209, 6.3743918644412, 
    4.37871328812049, 0.116417911321121, 4.45928928919066, 10.9862467275462, 
    3.13677075241324, 2.22535731533176, 3.91732272592089, -1.31066970187611, 
    1.44007358085818, 3.27786231467085, 7.90841452450894, 5.2698444425896, 
    -2.78748567398438,
  1.81034005932442, 7.3647873478557, -1.82206643802174, -0.152906185768634, 
    1.06473804920282, 3.08262556387458, 5.85950424855063, 3.04390727925414, 
    -3.14291001641695, 0.906695608579215, 1.36679317299437, 8.01247425667187, 
    -0.904590452111474, -3.14283612725588, 1.89034517682587, 
    2.53105954480284, 2.71940712842758, 6.20700733856788, 3.01345122191212, 
    -4.19155275829846, 2.57162682302478, 5.20603932868616, 4.79215567045332, 
    4.61540197097982, 2.22790154411362, -1.94758028729117, 1.64437909466381, 
    3.55672584317222, 7.33574842207417, -3.51221539797961, 0.920751216134061, 
    1.15971588542209, 2.86220726275618, 6.64448838963259, -0.646387406385727, 
    0.352465519788074,
  2.2870757681528, 3.53143685458529, 7.5555578096333, 3.30947506815018, 
    -1.07854424271512, 5.26612724023927, 9.53092183873845, 1.08955528019806, 
    3.85084931376337, 2.23389288241926, -2.21685714160085, 1.69979762213135, 
    3.32418343761372, 5.46141491346611, 1.64444130236381, -4.00516421301711, 
    1.67020294259317, 2.57752752807946, 5.60434717861278, 6.90954874168244, 
    -1.9370991081384, 0.478605961463377, 5.04490340594726, 4.82712666142561, 
    -2.54423775643694, 3.9633825566582, 8.96298225397022, 6.22281384825549, 
    1.08394314538844, -2.68264636642718, 2.95725777808116, 7.19195432308527, 
    5.07040263579934, 4.14085095718654, 1.45405982463088, -3.17163486293519,
  -2.41843121473823, 1.14931244262819, 2.2426557087436, 6.84947023114381, 
    2.07623630421372, -4.30656998059444, 0.456532316066405, 
    0.989708580367202, 8.34956213984632, 3.74287053291755, -3.53377474271306, 
    1.37740314294624, 0.323108704024854, 1.97063536239532, 7.6948566692801, 
    -0.409191411801138, -2.65726785427273, 0.37122358185251, 2.2368705337538, 
    9.79453495319599, -0.899694280503617, -1.2289727816108, 
    0.626119282733366, 7.55606832805448, 5.28126578505401, -2.78019628127056, 
    3.94338459831247, 2.03837768537374, 1.72039438356399, 3.3122381323806, 
    5.89097579175416, 0.899311946864875, -3.3506227996715, 2.33010804016319, 
    5.42587396011941, 5.38508748058851,
  1.12113629414632, 4.07210209148928, 8.7295489228134, -2.17362981206959, 
    2.05897698807755, 1.23584415806778, 2.47144705701544, 5.61391697951714, 
    4.33321595189527, -2.73122648011988, 1.11292607221109, 3.36427785955456, 
    8.46172503937994, -1.8048619665918, 1.48095913030665, 0.431355324927412, 
    2.21481115870115, 7.41342755079763, 4.42717829526239, -3.5478887568103, 
    2.55456061470974, 6.85559684061231, 4.31122974412742, -2.68916594412369, 
    0.751500621904137, 2.56348899351067, 9.25124846201203, -3.66478600383402, 
    -0.572664611511825, -1.10555342055106, 8.08472854521204, 
    1.81558197358358, -1.83156041488876, 1.85805187575609, 8.03447341159589, 
    -0.859421158658792,
  7.34318317566373, 4.79592586098132, 1.47123188934591, -3.61732514338445, 
    2.57614716437061, 2.48807843104765, 3.04351012856046, 8.50723318689759, 
    -2.27111248284965, -1.27944626285616, 2.0911202527494, 7.4281308729159, 
    2.49739902831152, 3.53799473190837, 5.08442787860024, -2.09830470906131, 
    -0.636411306609864, 1.19909434247572, 6.26425513522135, 3.99021307362256, 
    -4.18471635203399, -0.522662346606981, -0.642779338078983, 
    6.20145005148529, 9.72750931697843, 1.77417837498753, 5.27544653687611, 
    5.77580279316549, -2.01354466407921, 2.59700311890049, 2.00521397776974, 
    2.43588002337883, 5.08348274643276, 4.48915785543064, -1.08740832934021, 
    4.52091540115971,
  -1.53896696893807, 2.58797665861452, 10.5424925196994, -2.28370326685015, 
    -0.9289642610436, 0.0127014830018295, 6.67199229581268, 9.27031217253887, 
    -0.231765173729027, 3.63501858336591, 1.75745276192403, 
    -0.117034527410949, 2.97155595793948, 9.5648892690851, 
    -0.118988831225926, -0.493999516234146, 0.995345851493607, 
    2.1391099763271, 5.97942219930385, 7.35695297153259, -4.46750095509963, 
    1.95741628201038, 3.05351880560334, 6.49757067415584, -1.36423917265701, 
    0.69430480317575, -0.318543295406891, 8.63025085423353, 8.19014003863979, 
    -1.80318541741671, 6.39846223035559, -0.378809449161405, 
    2.17761315251423, 1.50849661198944, 5.81897838448991, 3.09293174985967,
  -1.62580522076662, 2.56148919851262, 7.0530874997732, 7.35736692179835, 
    0.343461578920575, -3.5809088288749, 0.856859031118597, 1.40453265581347, 
    4.57043606597564, 5.72037055756487, -2.3831463029414, 3.58893133892691, 
    4.37824193552106, 3.67907376725878, 4.89390519094474, 3.36415381586132, 
    -2.15737838371605, -0.548370209482471, 1.41274687956275, 
    7.99413186200313, 4.40509049127996, -3.27978665846959, 0.765664283645048, 
    4.9776486271631, 10.6461576435746, -2.13379905192431, 3.48382569078667, 
    4.34242261500154, 4.0657004851833, 5.55789779318547, 1.99798197456151, 
    -1.54629222014393, 3.52266192191216, 7.12303104975052, 3.8524121503263, 
    0.737726379483136,
  3.99975763191333, 8.80798365921629, 3.96140269144971, 0.0347872231669895, 
    -0.703374390218608, 2.21352115009014, 8.93206172537123, 5.66152806317264, 
    0.46652508814355, 5.39759287674635, 4.01389591510517, -2.41727405854971, 
    3.15045412863429, 2.72426249506731, 3.60635491812242, 7.51690597774566, 
    0.559538429325264, -3.0937096114232, 1.29395432337862, 2.36449042356371, 
    5.10027176072444, 5.28395165116342, -3.24541158089465, 4.55247036043733, 
    4.03555249378963, 5.06499246463194, 0.802302240296037, -2.1209928095093, 
    -0.923983232271687, 7.60098398289776, 6.12051002430397, 
    -0.99856955835889, 3.2916644445369, 8.65315227645343, 3.52342666790024, 
    -2.49909034299772,
  -3.51999840068106, 2.14234180860045, 3.87370478999673, 7.58009758121693, 
    0.0570347693974491, -2.958235011083, 2.91777092110229, 3.08507171276392, 
    3.0195200289818, 6.24177067876315, -3.38192342021847, 1.8878150692116, 
    0.0695833204346963, 2.99999095948135, 8.74474186479752, 1.61880308937782, 
    -1.35382234711925, 0.370837423370469, 3.03425319911476, 7.25705988165776, 
    0.653443944265528, -2.62435150927515, 2.08037058626098, 6.41228230671456, 
    6.29962866692029, -0.516030579521652, 0.0854678455659337, 
    4.41005324126955, 8.97200196907345, -1.58671895242095, 1.15932858610613, 
    0.454308130595617, 1.06964782843233, 2.81464043435515, 6.01127129356988, 
    0.976396536903961,
  1.77753682495209, -0.123703253934677, 3.44726299124959, 9.88001547616442, 
    -0.778919298642749, 0.808154888693017, 6.55986754650321, 
    6.29686119705569, -1.98488122420033, 4.90524443210488, 2.8610785739471, 
    2.40912611882899, 5.71892886867233, 5.64845000528345, -5.09757785921928, 
    1.34240867281122, 2.76450541162545, 4.13720374473599, 5.20403394418431, 
    5.35125530716597, -0.430382213136624, -2.143774041802, 
    0.0820942836889049, 1.61503998810275, 8.30814060771726, 
    0.377952693193332, -2.55978513688692, 0.46897068424894, 1.99101222210292, 
    8.22086107397245, -1.02826907144645, -2.26133750029398, 1.61749128723674, 
    10.3850862803317, 7.18994961838955, 2.20457736051925,
  1.79878385820989, -3.50473892494864, 2.11104224566903, 4.08279688911059, 
    5.77484400189637, 4.84768198979429, -3.14601759380751, -2.41725083448119, 
    -0.474841702125424, 7.93612600660828, 9.50302530458433, 2.9080805867115, 
    2.34716126220072, -1.33394660197943, -0.113123538564712, 
    3.62231139289945, 5.88739206272023, -0.810004578052755, 3.39883031235796, 
    8.72671600117095, 8.37054352808436, -0.208671537875754, 
    0.0713684633486249, 5.72769627620946, 10.5821026694556, 
    -1.12484573012268, 0.32365303531591, -0.118486732767289, 
    0.106240929842499, 1.41132988269582, 9.81744250937657, 1.84436665868131, 
    1.33839676616963, 3.81896263336283, 5.08324768824632, 5.73471114500652,
  -2.31203795377183, 1.67136299050971, 1.4077713427331, 3.00575620656311, 
    6.80856656684318, 1.75649920584106, -2.41214028380428, 3.68071688490218, 
    9.87590521937509, 3.29300566893206, -0.517625940164645, 1.62377288067773, 
    5.51119160441578, 2.70127990797807, -1.45486583692008, 2.93648841847992, 
    7.77468287669684, 1.72836547226761, -2.43246234456823, -1.29761749523068, 
    1.01526704179725, 7.3639388555407, 6.23324892641515, -1.24765285649726, 
    -0.0282798921582361, 3.13785066396196, 9.63515125235864, 
    -2.1216027976343, -1.46290333629696, 2.39316911144827, 6.06521494852255, 
    -0.952864893134461, 3.22267073952704, 5.50834618377539, 6.91853160131593, 
    3.05587037891299,
  -4.9472273567964, 1.31322192317452, 3.66680580581152, 4.70695876076936, 
    3.9236019912977, 4.7479473942167, 4.17093643773913, -2.74980523571099, 
    -2.91063224224733, -0.39012313015485, 6.3152941979311, 8.0062104895593, 
    -0.190084656090153, -1.77983195458913, -1.16654770462499, 
    -0.399393934730365, 8.25228677853021, 9.28871570304807, 1.42969219312968, 
    6.43303420378627, 3.43942956322981, -3.49453192622183, 4.11471848444804, 
    4.33533418537411, 1.90552835526071, 4.70821293468962, 7.39224150969534, 
    -5.51687127567905, 3.04331054130551, 3.17651824724061, 3.18823195930306, 
    5.12622583356294, 5.13965264468938, 4.01875471385213, 5.67076038999383, 
    1.75027087119648,
  6.62850856582441, 6.89866070791047, 7.03626401685268, 1.85329110308628, 
    -4.48127104655702, 0.189146548832924, 6.63960480586725, 2.46852388116518, 
    -1.54616301032026, 2.76288448341964, 11.1035380483175, 0.951152501745298, 
    -0.302744703059458, 0.537024451044149, -0.21973632222067, 
    1.85655493878373, 6.30465687990626, 5.67348010778391, -2.08217116421611, 
    -0.454633474206913, 3.10873063896962, 9.31274634903061, 
    -0.536692314793585, -1.36407840224876, -1.18059066243963, 
    1.92066268975471, 7.64940992809909, 6.06340821885424, 0.876012010210455, 
    0.131547810057005, 4.31054714198595, 8.02905864686877, 2.86556655033746, 
    -1.2318302173906, -1.73653469371157, 2.49903173679565,
  1.5068659698433, -1.87609665969385, 2.54943107787718, 3.80166245054305, 
    1.90223759593514, 3.92597686325512, 6.24396800012359, -4.43992693362344, 
    -0.234155660340021, 0.285831799001806, 2.10895069725169, 
    5.29621966880747, 2.94228724034794, -3.0164577745699, 2.34230581876353, 
    6.14508826248209, 7.1810774604943, 0.649047574910814, -2.28577703748264, 
    0.211944676868177, 0.15849889354746, 2.25335761348421, 8.39003083935699, 
    1.83288748826002, -3.64115602881201, 0.0451532626000244, 
    0.442055699245906, 4.49038979486023, 8.03168325854728, 2.65039001842808, 
    1.37295186841638, 0.51085457671649, -1.0423128919942, 2.43383824106742, 
    7.48301857940003, 7.7068680180311,
  3.04958062076139, 1.49621073300193, 5.95520928995119, 3.32402025947611, 
    3.34889387683239, 1.3279417942165, -0.841435553407115, 2.30753415298058, 
    7.14334213501904, 3.11762057759449, -4.40744434625158, -2.55159954521727, 
    -0.772965876227889, 3.25026322656278, 6.85596049584142, 6.63074417881829, 
    2.84433340358562, -0.479209881083793, 2.14246929777361, 6.79349071830404, 
    5.77550571796609, 1.22871150019103, 5.81391427191835, 7.85497162998115, 
    -4.83282527814808, 1.03027847014078, -1.27705956628068, 
    0.682634468649126, 4.63207281426313, 3.72985566758747, 4.27236102886384, 
    6.87379688943194, -2.15763584348645, 0.958365055750222, 3.90503730608699, 
    12.9386275922649,
  2.61045812772186, 6.92015185803606, 5.55343680094475, 3.12534903991089, 
    0.115972564583046, -1.79391427890097, 1.41019261149261, 3.5481714975382, 
    5.89995654443982, 1.5590748001163, -2.63628801692126, 1.86277634322209, 
    4.19318022959504, 5.71946718532722, -2.63596161333854, 1.17961634144466, 
    2.0884306193853, 6.72143691700928, -0.344346246250481, -2.97225497956926, 
    1.40063472267676, 1.91924786916632, 7.5187741252734, 4.08910572573772, 
    -3.28623899904929, 3.98944582810919, 2.99315265156791, 2.90156950214905, 
    6.40239119185171, 3.19698699329447, -1.98968495567945, 3.86272700624076, 
    7.89670872269965, 4.55164088329961, 0.485695496009312, -2.41142446066244,
  1.46280010445652, 7.52728166785324, 1.52349954623059, -2.9404302354617, 
    3.93538397590085, 3.24065028714407, 2.5774557050643, 6.6677777348754, 
    1.43873517035687, -4.80052916932007, 2.30602780907609, 3.63990964475763, 
    6.81755307361401, 0.469476833779606, 0.973235004866409, 2.46120855090933, 
    8.3254528000376, 1.87175204952544, 1.15193749611671, 5.42077981982918, 
    6.50683347764661, -1.56041571549667, 5.10804210052274, 5.13420113959599, 
    3.38591304799606, 7.11148233494744, 5.95617615750548, -1.56132862610277, 
    2.68284073553652, 2.24802061131236, 0.657566933217145, 3.0537558642886, 
    6.81108466178963, -0.820816691199934, -2.59878302175598, 1.37144910001386,
  3.99149238951517, 6.12957533126553, 5.97347352962602, 1.80297962855265, 
    -1.9285197840444, -0.66632192296186, 0.718109433612574, 2.94535223126365, 
    6.97967219051713, 0.597841170860025, -3.06380001970907, 1.30464079275696, 
    4.74816302700069, 6.94809790138221, -0.385616400133228, 4.89397017544861, 
    3.90670206979315, 2.76270047230913, 7.28003573385756, 0.0151967314265082, 
    -0.456493573501919, 2.04590825560134, 7.3847804240293, -1.03871097022051, 
    0.836383291513279, 2.33051435204528, 8.74222220010274, -1.21606391508672, 
    -1.05085509308125, 2.02025631267769, 1.86835446118742, 2.37917015652013, 
    6.65642402446169, -3.13252386690812, -2.44821140232576, 0.0924216076288369,
  -1.69247611597472, 0.876494480063388, 2.40592865204978, 8.19488928655484, 
    2.88897146414408, 0.360307713964445, 5.66069228508367, 9.13665637978161, 
    1.68953711028192, 3.66002835483419, 2.44616162940966, -1.2492797111294, 
    3.73093580420324, 5.78402819269173, 4.74073828218593, 4.42083202708249, 
    -2.20017982877342, 1.59769970439762, 2.76738389942681, 7.25545665093175, 
    -1.98582082903256, 1.57142315248939, 1.06123674881283, 7.4378785963253, 
    2.11540301570631, -3.95932941539258, 2.73348384388688, 2.0670519688671, 
    2.61250251390294, 7.68978891720443, 2.16348907021887, -2.90478159475444, 
    2.67667042922576, 9.19348960278048, 2.03190520999362, -3.20304470475557,
  1.30286981928153, 5.21192170668617, 8.80889942169403, -3.96134002815321, 
    3.2882730543406, 1.89865610714542, 2.19037411098092, 5.73024274684089, 
    5.71697910721194, -3.31973346474835, 0.525049130946971, 
    0.170209033640468, 1.37887897350073, 7.65250297884701, 3.44045965164438, 
    -3.3974113838661, 2.24093645861869, 1.56932441472744, 2.09755391796751, 
    5.25289285759507, 5.59408245766447, -3.71839527777149, 2.18207092537584, 
    2.12755111223515, 7.0293165228997, 6.23665058945678, -3.07908282546587, 
    3.56182042961027, 10.8294692699319, -2.49378898113739, 
    0.0914776982329197, 1.65831862596141, 1.25091416248925, 2.22157106617749, 
    8.29621571638111, 0.532339075428333,
  -2.41838275303687, -0.29374537266284, 1.47254644790221, 9.60237759241937, 
    0.52310537446921, -2.76665589050271, 0.611639707594655, 6.95340608392794, 
    9.25022918238226, -0.824254342105996, 3.24270042660137, 1.26581951390051, 
    -1.47788603765642, 0.430593547815216, 8.27961677527487, 
    -1.59212994711932, -1.56094992225531, 0.768659201210255, 3.7759957147218, 
    6.01143808000614, 2.32485840958738, -2.49559699466716, 0.885388425000872, 
    2.20346600323934, 8.53382009203577, -1.7406212279694, -2.31433423628184, 
    0.604803868191486, 2.67307532331349, 7.78138936830804, -1.66667568322837, 
    -2.04667007195341, 1.67065569282961, 6.33379740058621, 5.35354925199078, 
    1.4746536448451,
  -3.61840364011286, 1.63996689358257, 7.34790142443586, -0.501970223837738, 
    -0.617884018918645, 0.356932173126123, 8.34030279434768, 
    5.43346597578338, 2.65320294720767, 5.82578577843478, 1.58016356799457, 
    -2.16624287698603, 2.1768326857792, 6.76110577488359, 7.01829711142247, 
    -0.171389058032521, -0.0106070510845866, 4.92137310469598, 
    9.15272405827061, -2.11491968969508, 1.76193459462468, 3.73066018971509, 
    6.60695884387429, 2.12013853972986, 0.808700602964625, 4.99600389135409, 
    4.38805668985471, -4.05830441330251, 3.10298570287011, 3.26455516430819, 
    3.41686970947817, 8.31083847947855, 3.99244920244438, 0.651104335534043, 
    5.56749269607866, 3.94901851166036,
  6.86295050848909, 4.98069248196524, -1.93668153099712, 3.25070711793635, 
    7.73665823439919, 4.84930566029428, -1.45095134063002, -1.16693771423788, 
    -0.210284761311777, 1.80095445208903, 8.02446497854282, 
    -0.241472825546155, -2.15402676760101, 0.294915010190495, 
    3.29420325884652, 9.44677073550523, -1.40196531154366, 
    -0.315158873492647, 0.828989466808931, 1.38144366983124, 
    2.53163634202969, 7.57792201359897, -1.28029941656079, 0.846039920985757, 
    2.33572951276238, 5.9727791778684, 5.57466208541392, -1.01521040402774, 
    -1.95533361852798, 1.41435173553612, 3.59850262598156, 5.81019075716714, 
    0.947146337159738, -3.43686823760929, 2.18430936753436, 5.13220734857203,
  8.68929907651038, 0.381370678267785, -0.181160140362293, 3.23848662046347, 
    7.78458311119604, -1.55747241463818, 3.89116206281237, 4.67767061202168, 
    6.22191120451625, 5.73106924963602, -1.6387046855255, 4.41107746830191, 
    5.66060292511901, 3.85519615392443, 5.12596346301925, 2.42172019717252, 
    -2.87225481351312, 2.44495058796197, 6.46180996157366, 9.38368547360647, 
    0.435913395669178, 1.68341075653663, 5.34247747419023, 6.65750543340941, 
    2.30026976151659, -0.856436207320341, 0.210058157827784, 
    3.10684308322256, 8.90209106870202, -3.55059144800686, 
    -0.195101413283781, 0.0420639880441311, 7.63008250699018, 
    -0.0334508458434581, -1.14109972624408, 0.422313360707202,
  -2.27902293048076, 0.948895688580944, 3.88909431438193, 8.35392679368212, 
    6.14225076939671, -0.0122935463618985, 5.96462660500357, 8.1652139756392, 
    -3.10186695455229, 4.04557284484244, 2.8265998414494, 1.96043740789591, 
    5.56948948371795, 8.15168912113404, -2.00952885357694, 1.53108017256553, 
    1.86783860057332, 1.5176120525834, 3.29305432584998, 6.40740769536053, 
    -0.00274891885055739, -2.20338464821297, 1.36419742886449, 
    4.43258408394694, 5.77240502391391, -2.45128640562552, 
    -0.477985119669136, 1.09554486075786, 5.06599993169851, 5.26541240666641, 
    -2.8251750244811, -0.450627844428047, 0.916877608142568, 
    3.26032878450197, 6.79580202432135, -3.29378038277066,
  -1.92674869591138, -0.463346702083165, 0.578263950542125, 1.4317277231195, 
    2.97045221856487, 5.65624162055293, 0.123327923766473, -4.24384428379246, 
    3.53837084839724, 3.26279939672967, 4.17007960826365, 11.4772375116724, 
    -1.21382012053809, 0.472642074920477, 3.46812951473731, 5.19565916092251, 
    4.85279412784151, 2.20658581834661, 2.09052749610643, 4.98987217581831, 
    3.62243520650105, -1.81706517562933, 3.46404722625011, 6.56518766232849, 
    5.36182020453928, 2.34452708185294, -3.1600250772861, 1.12163398515499, 
    1.03336491786512, 11.0090225067091, 0.948219946802737, 
    -0.486739862230353, 2.60857934734444, 3.4909043062376, 5.39054756791273, 
    6.33127953813601,
  6.26031142078113, 2.51056862921971, -3.25839083202483, 0.11660204677397, 
    8.92104651220262, -1.61756301270476, -1.45355331850669, 
    -0.0988308329414487, 1.75974418530892, 6.64167556995426, 
    5.78459930143459, -1.71205165692681, -0.562655486912453, 
    -0.424856361875109, 1.4614736292328, 5.16047743410244, 8.45976766574992, 
    -0.578764510177014, 2.50624508806366, 3.89468166240965, 6.10951342337614, 
    5.12316093688303, 0.686768928648661, 4.47163670174982, 9.42271445371146, 
    -0.105422235364814, 2.34163578500919, 5.74250913122151, 1.73358153748028, 
    -1.31266419411928, 2.39727547522567, 2.98824457641522, 6.04258545066748, 
    0.130892894608692, -1.57667197742426, -1.7074107249772,
  3.57714676752179, 3.25888725762195, 2.87121381548036, 5.99023307928986, 
    4.59546350753946, -0.177158470038949, 3.98922502077442, 6.67059000380388, 
    -4.38786566343663, 1.22275552790085, 0.471929967619101, 7.2700505799637, 
    2.99585015639792, -4.46476714456226, 1.84159094519486, 1.06867725546874, 
    2.04654640007467, 6.26773401590725, 1.62955657982134, -3.3050118253676, 
    1.09286661453937, 3.74768023588432, 9.18745253246596, -3.8202115564069, 
    -1.3541116511959, -0.901778453360451, 4.88166926492758, 13.4256061341288, 
    1.09849424836302, -2.29174423116242, 0.468695140854241, 
    -1.18633988641508, 0.117682617372691, 6.24149913102422, 9.08886166343665, 
    1.74691266933281,
  8.42841061668962, 1.66997709547302, 1.91938665579796, 0.0860724037368397, 
    1.50970324362431, 2.82278412081828, 9.80462442130777, 1.17842285630483, 
    -1.99426040946628, 4.5414383013748, 7.66294547809637, -2.12143509952526, 
    2.12785860050094, 0.83472983979398, 2.11643027856518, 6.37017883313064, 
    2.7581526106179, -4.43429681618865, 2.32601698010928, 4.02660619009605, 
    5.02679040090592, 5.70845096463642, 1.02228422992767, -3.10014428026647, 
    2.18069823410402, 6.42355358717717, 6.92521379984502, -2.00869250138332, 
    2.63521812368386, 2.39613585129038, 4.71954960681726, 9.44815725292673, 
    -2.25593501259069, -4.90750630660573, -0.689024194165835, 5.2589244730759,
  3.1127494562016, 7.44793250893171, -0.730955677557605, -4.42065967353707, 
    1.49713033856176, 2.93893687341075, 8.4940739581825, 5.38765012899741, 
    -1.16030472561288, 5.37115142084264, 6.92282152714977, 3.49281559944802, 
    6.05245329602301, 2.63344804428799, -2.61851073613908, 4.2135018216353, 
    5.67035286734995, 4.49355154389611, 4.89077335737145, -2.20079472197139, 
    -1.79766442325884, 0.390396067977409, 0.546228646398831, 
    6.14062692456063, 9.47538109694205, -0.737055972033423, 2.36559507825878, 
    0.354086725505665, -0.369879262864405, 1.28041132771609, 
    4.87031529670441, 7.82431432193154, -3.73888946921622, 0.419823862510739, 
    3.49266624817635, 2.50877776385285,
  2.44596232263325, 4.96062695347969, 5.15674952496275, -2.82417662836753, 
    2.88084903862502, 3.57588935822987, 4.87795361927742, 5.51050705697752, 
    -2.3784778249592, -0.785326275299367, 0.34533565371333, 10.9971017654633, 
    1.8748758521082, -2.20419978726381, 2.26556508366202, 0.769368696553068, 
    1.99958835337991, 7.26101447687406, 5.8333406412572, -0.199387386192685, 
    5.14558509454003, 9.52971651151683, -0.395263368267275, 
    -1.11549440132246, -1.19217091747444, 1.46668586874125, 9.36922182076079, 
    2.83849301802507, -2.87149687766781, 0.604518620031941, 1.00716118901667, 
    4.633658366197, 8.50020636285963, -1.9689594591641, 1.21920899984455, 
    1.5630763539358,
  -2.09812741855334, -1.79326576662454, 0.302037054565311, 0.527597831397547, 
    8.44324322840809, 0.616169901230633, -6.47965072283797, 
    0.799121885023505, 4.77023872498772, 10.2258243337356, 
    -0.0651804343169382, 0.477863108622435, 4.83109831728968, 
    6.17529516452062, -1.4411898768487, -0.51917217346246, 0.760836058742869, 
    2.88843142702254, 6.72887095534761, 2.89804852816655, -3.07813879265411, 
    -0.273247446156175, 0.717869298840538, 3.06407104444151, 
    7.31957769067805, -0.0372011053941215, -3.791576901639, 0.84720376434085, 
    4.19130101662165, 10.1433704205172, -0.511073504841812, 
    -0.536428427697294, 2.61717939889795, 1.55480605731398, 3.36503431875742, 
    6.47512768207641,
  2.1367203610352, 3.51921382157307, 1.33026372880308, -1.05481390923727, 
    2.77359762551224, 8.27100694128882, 3.99060952964922, -2.43990590243397, 
    -1.67404014624149, 2.69738599289792, 6.37452586913952, 5.4397570168431, 
    3.67508224714181, -2.80969476839374, -0.0266689044738646, 
    1.11066736658677, 10.5709654111384, 1.36388518581069, -1.42999138265325, 
    2.31064643413034, 1.5896936442893, 2.97372628230207, 5.84320501461178, 
    -1.17869976151253, -3.797938389562, 0.936929336491391, 6.66343572672763, 
    8.76482552468434, 4.53194153731408, -3.7311529510712, -2.7247193670914, 
    1.20513748886757, 6.75381712350097, 5.35632139496523, 5.24340435088132, 
    5.00032789010108,
  8.90353261075169, -0.736210515298732, -2.93142557588034, 
    -0.731681653346076, -1.45578072664995, 5.21080279422145, 
    8.21472460160208, 0.829003554664283, 5.00042713006163, 3.55151164426379, 
    -1.5682852772518, 4.49332649799021, 8.09174469750894, 4.57123938664108, 
    3.6534620780425, -1.33954855917123, -0.898251394247768, 1.57929026365409, 
    3.83062132737761, 6.72085120618902, 2.85407209890563, -4.86631007135235, 
    3.4221849918956, 6.0131801761213, 6.36776599987141, 1.61589947093979, 
    1.69944937606523, 5.43956515255214, 4.60244867818777, -0.95313117602243, 
    3.54270311467865, 7.65358504689767, 2.38388099533316, -2.32555660353349, 
    -0.834170847318072, 1.50955308168613,
  2.40574342897687, 2.92060970699947, -1.06620687208278, 2.02176549371466, 
    6.89281767403183, 4.94239345318678, -4.38325668350109, 1.94400231153085, 
    0.804262356127675, 2.51660626493755, 6.68092737877866, 1.49822469567609, 
    -2.79012253271785, 1.79961991383403, 5.55226910523616, 8.04709730185963, 
    -2.03417839570903, 3.01110003120032, 3.58323493643992, 4.9020959777099, 
    5.97079632222635, -0.370541345472847, -0.683091063869835, 
    2.61248016693234, 7.3172454650878, -3.7814347120587, 1.90534573296872, 
    1.93242748503459, 7.38791404992629, 6.1216204530506, -2.85214951915675, 
    -0.627945352172281, -0.583685144252841, 2.46264119507366, 
    8.59823929999283, 3.69413025640675,
  6.38613261672377, -2.34047712861021, 3.8025936506916, 3.99116156086044, 
    3.70536786167403, 5.75524455102049, 2.72236032506713, -4.14283517494362, 
    1.7643957017382, 5.84728639478418, 7.9901768645315, 3.08258689417461, 
    0.646311920979246, -0.21067147197784, -1.18793505910195, 
    1.61337060420996, 5.545979036778, 6.36411997225568, -1.2290847842022, 
    1.53019574290168, 4.76853643441127, 8.71693257069316, 4.14639647954409, 
    4.43945399174298, 4.28169268049763, -4.07600045421273, 0.969425667797881, 
    0.425118263515371, 0.68179379681812, 5.67997567226647, 8.20364579780824, 
    -0.80166743321141, 5.04374900528184, 5.08401213599003, 1.01373633155223, 
    3.73696878570162,
  10.0096999777338, -1.93651898791297, 2.22526039282129, 2.6743738272383, 
    3.35237196550146, 6.54132943817133, 4.28000145292951, -1.80389117101268, 
    4.40589704688493, 10.5812254103754, 0.384597477684614, -2.11367848194909, 
    -0.595669225818118, 3.63788787125774, 10.0036520618832, 2.40702864896624, 
    1.90539992860481, 1.69003565051078, 0.242910074396303, 3.31064266440729, 
    9.09516125793343, -1.84328131728922, -1.31498633403245, 
    -0.0312054802430852, 1.66770416177607, 4.08501896275306, 
    5.81273731360123, 3.91697794830758, -1.37690279883555, -1.23415906815034, 
    2.88320209293989, 10.0891848391245, 4.149587178347, -0.895385738753437, 
    0.637762782916503, 5.55242159329311,
  0.727238275761411, 2.97491457012678, 6.53818840013148, -0.357092413353175, 
    -2.91271586515828, 2.13994970002549, 7.92462498686508, 5.44238092914199, 
    -2.40006200467868, -5.26325674913769, 0.729164196803663, 
    5.68025984273162, 6.89328597006551, 5.67042068422348, 4.14199596656717, 
    1.8292222345716, 2.15855218553893, 5.36701274794071, 3.20617300702808, 
    -0.270894431610755, 3.35825816208714, 9.33810048812912, -2.827934949521, 
    0.694085821542878, 2.96041659041742, 2.44737561966355, 0.758827331987435, 
    2.20378048521349, 6.97022489094691, -0.69492112329394, -4.47389579402469, 
    1.24765724859537, 3.99562579895487, 6.1044050824364, 3.26193848969216, 
    -2.29470035853251,
  3.46264993109954, 4.47702411945699, -0.297705134002423, 3.18623691347131, 
    5.96256637109051, 7.30786348576393, -0.822399598503596, 
    0.422788043128548, 4.18608594084814, 9.6309634925402, 0.39522496733591, 
    3.32561147715162, 6.48811684406339, -1.62319399849812, 0.953281827925774, 
    3.10191364658877, 8.34448905858251, -1.6410124739617, 2.40381950861709, 
    -0.186424917121988, 0.808025301924348, 6.53434479503378, 
    3.02113911345021, -2.7186597635029, 1.93693918960881, 7.45940945077367, 
    6.36084387421763, -2.16876323452919, 4.1338969312088, 7.84236996641494, 
    -0.126590250933226, -4.82228495132982, 0.467439490845778, 
    3.11586780158423, 7.07539742055679, 3.58818656238643,
  6.25157341821806, -4.03630886820087, 2.95737416139436, 1.88240347986782, 
    1.46683817924306, 3.20170144622056, 6.26773407567077, 1.05756780711328, 
    -1.72301114466957, 2.50755194861739, 7.4100233847818, 0.0306836472962868, 
    -2.60459598469452, 0.530580022191915, 1.52939067473276, 6.79395070782524, 
    1.32786778738056, -3.78936164801798, 1.72782061872408, 2.61827398994715, 
    7.13076276724773, 4.13102599146301, -2.54338073631024, 4.34978035986867, 
    8.79041104448964, 3.30655172250494, 2.89885883393794, 0.751894752291939, 
    -1.57452472659363, 1.97423472782882, 7.86251064614851, 3.48469590306333, 
    -3.859548088896, -1.64205570475058, -1.25233344212954, 8.32031442520611,
  10.2051188151957, -0.599623152998424, -2.69776484510563, 0.373618129703898, 
    0.104847206622596, 3.37832769914368, 8.22755453969931, 6.02050618416207, 
    5.48560639722944, 5.41884702702384, -0.250616232262282, 2.7256702352791, 
    4.29347180456558, -1.90308158323498, 1.14176123094863, 1.18235629578159, 
    3.37273392829533, 7.81612455139198, -4.84164964247705, -1.97778453643119, 
    1.15347503557963, 3.4226046197743, 4.3951826664011, 7.47317892645715, 
    6.68429407431258, 1.20019718876044, 1.69986411583563, 4.42336587796036, 
    4.04833970865544, 2.35185626733525, 5.71123126693196, 6.16215939800854, 
    -4.75795272172012, 1.48457264588238, 0.159845867094476, 2.86690118727292,
  -0.940397130278678, 3.11050707987498, 5.11537410601504, -0.416089785974985, 
    2.30047431522131, 6.77977372188564, 5.82190522738419, -0.963190597999186, 
    4.59214820262736, 8.59162388814616, 4.07521908357781, -0.541504082382714, 
    -1.74542790982242, 3.01579521920714, 6.96951087184915, 4.42549691478196, 
    3.35786740915388, 0.942180750237231, -1.6974983417853, 1.52695388295482, 
    4.02510072205513, 6.35123390704078, -0.505292336429553, 
    -2.65757624598058, 0.924551651752636, 3.24893694680266, 6.9165343081584, 
    -1.51515756429159, -1.39616331192109, 1.1250697139326, 8.01186317501762, 
    4.03704892936773, -3.37811016041128, 2.33638519042852, 8.59218316795796, 
    7.73428574231185 ;

 Y =
  0.00204997293723586, -0.0497989321436717, 0.0291962363495011, 
    -0.0131350303202905, 0.0203595329892491, -0.0390429888075219, 
    0.00303253064020953, 0.0195957852700742, 0.0150166113192463, 
    -0.0375352351217682, -0.028194794400409, -0.0561420846010276, 
    0.20377076197604, 0.445637947032072, 0.134744286883157, 
    -0.208936102609338, 0.240260418275767, 0.491499090863347, 
    -0.238096214568055, 0.138412364481361, 0.752392529461686, 
    0.268194494105024, 0.20299071299184, -0.0194163274582493, 
    0.703654254313394, 0.594954521129343, -0.552849494060506, 
    0.128297271248023, 1.04132142550953, -0.00413747932087959, 
    -0.104186221509653, 0.136843740334649, -0.167244791689055, 
    0.125267013650451, 0.0798416065272884, -0.0203316794011367, 
    -0.126441367401794, 0.00273161683052997, 0.110227833611516, 
    -0.191646136936242, -0.103102150540925, -0.0958733770148624, 
    -0.0302550531302221, -0.0833919423301146, -0.0296798856221585, 
    -0.19094567280079, 0.015368367819517, -0.170772329486118, 
    -0.0333350267538376, -0.157234404158521, 0.0425154916899873, 
    0.0275120668238928, 0.0591880062536501, 0.0160108885455187, 
    0.0419982261814824, 0.0169846481375218, 0.00815398500977522, 
    0.033165226572601, 0.0221782256891696, -0.0121206572821519, 
    0.0594992311776675, 0.0911944895899721, 0.0995283439743617, 
    0.0841530127080123, 0.102271302665816, 0.112254743731293, 
    0.0663964382667706, 0.0444038221667676, 0.159454403877659, 
    0.10790953640384, 0.00278024860072358, 0.25406899464573, 0.5458115502716, 
    0.141533143152305, -0.22519511297407, 0.50139225488943, 0.55481011739886, 
    0.263586545358839, 0.195770178473097, 0.611988840365391, 
    0.331701450051767, -0.456963409867098, 0.271893307474603, 
    0.585661805308727, 0.120744495747801, -0.272415597830285, 
    0.576424397597834, 0.956662529020158, 0.220959369055226, 
    -0.0381105138036277, 0.0244216708817248, 0.129577385102126, 
    -0.0609845177849229, -0.0649828896946118, -0.0602116936848863, 
    -0.0922503739760802, -0.0584834549748304, -0.0212251775033779, 
    0.00188787483392186, -0.210977466991514, 0.0962174704823078, 
    0.262468552488366, 0.203588409054107, 0.10080646010215, 
    0.0076370182391855, -0.028275664970401, 0.194790308537264, 
    0.367962120500715, 0.292825816277693, 0.146712240506941, 
    0.0214100389304712, 0.135745839241113, 0.199679723165341, 
    0.192349313574468, 0.175557776560615, 0.0945126723764671, 
    0.105843255580183, 0.306307136174986, 0.285101685095638, 
    0.123400915071458, 0.00915930277432729, 0.0653236466341563, 
    -0.0603711536264322, 0.0478764054077974, -0.0144327836911175, 
    0.0543027971642698, -0.139731361616028, 0.0140624451884662, 
    -0.0812827635316473, -0.0979191427057691, 0.0467217105044994, 
    0.117841554302519, 0.040033306659669, 0.0429069501458206, 
    0.351686361228346, 0.188823582160906, 0.0577470544101083, 
    0.399914338493784, 0.0602641101780935, -0.0359149663786647, 
    -0.366639483645313, -0.0131888965057228, 0.838567775757481, 
    0.0352458840257181, -0.432205767077031, -0.130131266016592, 
    0.849227311576768, 0.168454754203689, -0.241000788474583, 
    0.399381675217721, 0.57821057253061, -0.125452902682838, 
    -0.149186001018304, -0.0767801630085281, 0.394893831548943, 
    0.0171977488489317, -0.118279372782205, 0.261153309548124, 
    0.0126987814111994, -0.0737090490933939, 0.0481286072244767, 
    -0.215967855137001, 0.0943068637486173, -0.255019955689472, 
    0.0417476619881787, -0.320152799016366, -0.0128225622325063, 
    -0.23454649762644, -0.0162499965560928, -0.231100094250533, 
    -0.0246778940779629, 0.0550389806685299, 0.0465935936279484, 
    0.0579565396745373, 0.0732921723421118, 0.0764312273959734, 
    -0.0205271387168536, 0.119847911936448, 0.106821308975725, 
    -0.0373933159343649, 0.0988337930588616, -0.135035474018321, 
    0.314391336559378, 0.313595466584319, 0.294593182224817, 
    0.60782062493324, 0.342409380342032, 0.0880308488734187, 
    0.0281514547896345, -0.0797236271485396, -0.482532757154356, 
    0.101498250909603, 0.913059767065751, 0.4085102768377, 
    -0.124873179897668, 0.831553971215362, 0.492763960819414, 
    0.534129855109847, 0.933964491891264, 0.205458494847947, 
    -0.0853684514860638, 0.0212924521795493, -0.00880275700731657, 
    -0.00271244797585451, -0.00385803556405623, 0.00260084937283328, 
    -0.0216144648137182, 0.0851766777104446, 0.170343036962807, 
    -0.166552355839782, 0.0914685694800735, 0.392297732822024, 
    0.200511101834297, 0.0565296363578558, -0.0548598038000972, 
    -0.14649786770879, 0.15809676863057, 0.486259378100235, 
    0.433830761919926, 0.124733045373979, -0.188381080455926, 
    0.0134835075853222, 0.477238520550528, 0.128322436498025, 
    -0.145833156118023, 0.194819179260448, 0.345701457997333, 
    0.0906699195594333, 0.0881055857296815, 0.441422080297968, 
    0.199635682487993, 0.0746191127510022, 0.045713761217047, 
    0.0442700076140147, 0.0489978097580561, 0.0494439601607399, 
    0.0478739744261932, 0.0563571094421352, 0.0411952703717918, 
    0.0173537078521519, 0.129734758620474, 0.0443414755336963, 
    0.0901866108502833, 0.362925836779857, 0.183303312749551, 
    -0.013834003049639, 0.0960015878342071, 0.345683578478068, 
    0.127888971507709, 0.314202432356724, 0.38518832866643, 
    -0.110069764194775, 0.0609203484968263, 0.416757388707711, 
    0.602979136780169, 0.348989283598245, -0.08257035568209, 
    0.64001047729377, 0.267026003703362, -0.108974450498436, 
    -0.25461456037015, -0.151603463257085, 0.0294248280859118, 
    -0.247233396967888, 0.0108139967569543, -0.235025851119094, 
    -0.0973991460549526, -0.123185242051234, -0.00555820348756006, 
    -0.194789068265301, 0.0786683101879924, 0.0815161149041453, 
    0.15754810545673, 0.16996829871166, 0.178015776154407, 0.197829402859416, 
    0.172109444887568, 0.22438353539426, 0.19933847966714, 
    0.0929903498478263, 0.0308022892831271, -0.0158178726991642, 
    0.0452901414185048, 0.030964172804951, 0.0136514171402696, 
    0.039221733533225, 0.0724012350890243, 0.112496218729943, 
    0.0658154285244752, 0.198308313031424, 0.0611627044354236, 
    -0.207109115752705, -0.236337704962647, 0.752937076444948, 
    0.318469272073788, 0.0397480076643001, -0.255561451548192, 
    0.115701256728128, 0.535437724337542, 0.438199967957117, 
    0.263073372773402, 0.163268248450016, -0.0292922698349016, 
    0.252001163902626, 0.312378924292924, 0.063476578572174, 
    -0.121622351030963, 0.199675940005847, 0.368627399254184, 
    0.125917129307319, 0.0311415385711861, 0.0332361051004112, 
    -0.335937120709526, -0.0247228314455235, -0.253739020482159, 
    -0.304675087458347, 0.0831070297727441, -0.0925484900402814, 
    0.0816298669851626, -0.316465850615294, -0.0159842706214783, 
    0.0480264886085068, 0.0471429150900659, 0.166101468820899, 
    0.181528465220068, 0.0515560284700833, 0.0756651293917344, 
    0.356661777784697, 0.130947274540358, 0.013779340135619, 
    -0.058239852037008, 0.403368811764161, 0.234398679988001, 
    0.0887300767962117, 0.804980608357893, 0.374112988066207, 
    -0.150930312489169, 0.501390366257005, 0.706262330475588, 
    0.186496022859161, -0.10986350046044, 0.276962730834899, 
    0.744967864517137, 0.21345421683307, -0.285938477865857, 
    0.217822669588111, 0.466205924471136, 0.149861345255454, 
    0.0245758848888921, 0.262851630565369, 0.364798209523292, 
    0.275133622440131, 0.0910601332160764, 0.0438207322392835, 
    0.221373308563667, 0.0172360725966095, -0.0597269746558063, 
    0.0245462701926907, 0.144029036041253, -0.0412384938092435,
  0.597235175577898, 0.377443757897011, -0.249236699433216, 
    0.572577543360787, 0.844988552617347, 0.36730937467186, 
    -0.153977346448673, 1.03847075912008, 0.396515541223608, 
    -0.0366049952034842, -0.244676020790342, -0.256731214323015, 
    -0.0288058246419793, -0.27052203242509, -0.0637333241639248, 
    -0.277488240552575, -0.038122309292852, -0.288349451965718, 
    -0.00963291743000244, -0.184372469267673, 0.192354888490774, 
    -0.0799915090007096, 0.101085768433791, -0.137562362338435, 
    -0.0196322217121049, -0.167208243836931, -0.0825237149388971, 
    -0.0341040895072051, 0.0740212550460232, -0.180036770996569, 
    0.0572526556727272, 0.0613454495557156, 0.063851919350396, 
    0.0880833064901165, 0.0752130786990197, 0.0786893649007212, 
    0.0663631362293113, 0.065730419302772, 0.0813333968788909, 
    0.0774897030621383, 0.133313715145163, 0.147227614487929, 
    0.118504760960606, 0.116808432596785, 0.115186058983971, 
    0.113903489987224, 0.112657365973707, 0.131343820095705, 
    0.118367268703868, 0.0771978991131493, 0.114438661904481, 
    0.140570269908696, 0.148391419117489, 0.192983374245029, 
    0.204548184616529, 0.154819352437992, 0.183886491647629, 
    0.223626222865467, 0.152315809616634, 0.349470014856258, 
    0.333012221934986, -0.104819232570803, 0.231678128646268, 
    0.658135136889408, 0.0889912794013664, 0.107233682731343, 
    -0.239515065026216, 0.0237340176898688, 0.535157913025918, 
    0.301753928501181, 0.21538276740006, -0.415695306275495, 
    0.491263071311345, 0.395277414639777, 0.0483446415139575, 
    -0.220519069002675, 0.240626064070234, 0.576848104488295, 
    0.501446945798132, 0.329084305123641, 0.135859458899245, 
    0.292653976300353, 0.192567287627909, 0.012910804088538, 
    -0.0238079652256599, -0.0531881012142569, -0.0155811226376939, 
    0.0316513335218746, -0.01023436638936, -0.0598177059924049, 
    0.0280353672267552, 0.112919115215591, 0.147085663038067, 
    0.184075649735922, 0.185510162903347, 0.0564995810557861, 
    0.194101337737398, 0.451209610388453, -0.00314374159656031, 
    -0.0350504929733749, -0.285482163349303, 0.231906415523501, 
    0.475692391596928, 0.361945649551793, 0.20960745834247, 
    0.0452423546566639, 0.511703523788789, 0.220148338590597, 
    -0.0534645635074312, 0.0820094841539807, 0.347358476715145, 
    0.791231630370502, 0.450875484664056, 0.0942662259390675, 
    0.127383554035854, 0.199015406571853, -0.0478649773001324, 
    0.121701482760676, 0.187669039341443, -0.0599978709886112, 
    -0.0183447516297674, -0.268148403072631, 0.175915602356718, 
    -0.15127799152674, 0.105106537038949, -0.257631998248972, 
    0.0724288548516835, -0.124874780951011, 0.113181300878254, 
    -0.370691879611799, 0.0389084864891939, -0.0366348524173652, 
    0.106423940086837, 0.130955947236774, -0.0389567485023394, 
    0.0535898077923081, 0.302216544516032, -0.00825322085103598, 
    -0.0392620322109448, 0.0244105628317148, 0.275939050353662, 
    -0.393688299312165, 0.0895888752099895, 0.572814826274225, 
    0.387173780542817, 0.31290648197123, 0.278427144872743, 
    0.0958485372841915, -0.482807823461263, 0.188028471956841, 
    0.530996437928736, 0.338055924029098, 0.506513292116053, 
    0.341553457794838, -0.193564356890207, 0.0396017555049353, 
    0.689527927314345, 0.0974915755993024, 0.0372347619223951, 
    0.0194165038586265, 0.302500709603573, 0.176561742257021, 
    0.102014807597462, 0.0852509775513179, 0.176490162952726, 
    -0.0659885282376522, -0.0134251209587467, 0.29232653942564, 
    0.3189361997959, 0.122955352165942, -0.0212860892587077, 
    0.078378544498503, 0.29051559196816, 0.070921817937083, 
    0.368493651088373, 0.446261039464313, 0.0063625558919235, 
    0.343909869688884, 0.639229960271526, -0.00756060219617177, 
    -0.0715133188596028, -0.0210681920641239, -0.0326843076740113, 
    0.0282738410393625, -0.0590402079123725, -0.0751213139877788, 
    -0.0090521199719668, 0.0284671352654538, -0.0886928577874761, 
    -0.0456695301074078, 0.0335128828195841, -0.0595963227314362, 
    0.0399363845545203, -0.0134140173198846, 0.0416889531012339, 
    -0.0376027909318482, 0.0261638500000899, 0.0296936973148744, 
    0.0852488660582239, -0.0858403798013574, 0.0898066834085362, 
    0.155073629253256, 0.0648600968607886, -0.0215338194373529, 
    0.1505891300714, 0.359337558483065, 0.118841222488518, 0.114213643540837, 
    0.321813816524512, -0.403222776442922, 0.560515115487967, 
    0.449342443025994, -0.147733433453776, 0.160968197086115, 
    0.782911599011634, 0.0496487350222884, -0.258409862786077, 
    0.262795481340242, 0.616617246383456, -0.131456175110291, 
    0.0632061166510069, -0.256410395954445, 0.34423961247549, 
    0.0338142450618976, 0.0804757390717396, 0.153214988481417, 
    -0.161775693794341, 0.150249877372137, -0.059539412326204, 
    -0.295735928399206, -0.104163543175198, -0.173393600707523, 
    -0.0416616423402965, -0.167751749784901, 0.0659192843942806, 
    -0.203743471846298, 0.0719318041799099, -0.147085674652452, 
    0.0470688456265986, -0.187777984028049, -0.00111220958972019, 
    0.0453156604399614, 0.0619501352842376, 0.0614068348443555, 
    0.0699743377212849, 0.0619075849474553, 0.0538046966863108, 
    0.0557648807573963, -0.0457136055563601, 0.095700909413056, 
    0.37199055212679, 0.0668453605932305, -0.20294971022596, 
    -0.00422820720414474, 0.552323913764524, 0.201833268814015, 
    0.0689204691668964, -0.159403003121724, -0.0204205469787287, 
    0.63311048457113, 0.0838470180663057, -0.0533148142308137, 
    -0.396865303767326, 0.0658158421818265, 0.544401872262784, 
    0.437822255654542, 0.126813332105667, -0.400218711798309, 
    0.0265199627444057, 0.415977357089761, 0.0580986978156717, 
    0.0560731627569898, -0.0549354107176556, 0.115463802970391, 
    -0.118863732745161, 0.0822894799738095, -0.472062675786815, 
    -0.0749169134341807, -0.163105724416494, -0.229636012864629, 
    -0.0115333633341319, 0.0968871472202706, 0.153989516516116, 
    0.204969536128761, 0.294226277907041, 0.303450428240275, 
    0.205591378860499, 0.14557593014766, 0.296819457759756, 
    0.366295387086002, 0.244560703075844, 0.17626697123723, 
    0.158383050692896, 0.167673207797787, 0.172499382578893, 
    0.140384307618968, 0.133442354696348, 0.170117620040467, 
    0.177291399033447, 0.134190801006693, 0.129481241021742, 
    0.136627377053132, 0.1062070467559, 0.173178655833523, 0.250488093629332, 
    0.152081989832996, 0.0478599387822261, 0.17270024118602, 
    0.286820056320493, 0.29424775520509, 0.165478578599543, 
    -0.113181904698563, -0.0463986910922653, 0.465605446865572, 
    0.268932121682236, 0.149529842134543, 0.123987792931919, 
    -0.241641835385926, 0.139152164802306, 0.452338370507446, 
    0.332190868263794, 0.169772307939928, -0.114930739864295, 
    0.121606709720224, 0.191543887503795, 0.373627693399468, 
    0.288350488905698, 0.231207081740644, 0.330457415061758, 
    -0.169649283942893, -0.343639974546677, -0.0762164806906365, 
    -0.196502689260745, -0.157426641645007, -0.156484526855873, 
    -0.159825853284811, -0.106618076071133, -0.165773737222848, 
    0.0123564471164707, -0.195225381832063, 0.0685067114969654, 
    0.0372643709972608, 0.0556930954875858, 0.0707898426987124, 
    0.081095831040307, 0.0519321889526801, 0.0781920989788919, 
    0.0722464822919294, 0.0653708684100384, 0.0196345712848705, 
    0.0154150388674709, 0.106495360388596, 0.198475938701148, 
    0.132963273060647, 0.0314725104518938, 0.175627419797484, 
    0.161610660862324, 0.267759201311189, 0.347752059170986, 
    -0.180845868670765,
  0.459866265285988, -0.0940249697150692, -0.0891346838741359, 
    -2.55739868842142e-05, 1.16343142656354, 0.800409991888862, 
    0.155887366047107, 0.770575623921884, 1.13523439105425, 
    0.310011501442104, -0.108814293632201, -0.28160498623039, 
    0.105253455068834, 0.0142137655223242, -0.147826579347833, 
    0.216298472227029, -0.135347286736392, -0.206978357995283, 
    -0.234343409713677, -0.170278801237641, -0.190746490027716, 
    -0.0994723186406062, -0.148452043353491, -0.174228865827452, 
    -0.0133370846777774, -0.166117376740666, -0.00612873633274962, 
    0.00802560367717677, 0.11065179555369, -0.238242905896009, 
    -0.0350987358954939, 0.264626933838818, 0.0026808780443992, 
    0.095934734117988, 0.336330000423913, 0.161821682118438, 
    0.135657397818668, 0.358402225072555, 0.0148786155217161, 
    -0.200608459495732, -0.239377105732539, 0.203462430014633, 
    0.594087111376117, 0.613165514993532, 0.309367312867227, 
    -0.046491991253832, 0.790803525276923, 0.627434545793895, 
    0.114908934628114, -0.102096890151803, -0.202731571621029, 
    0.421781702800318, 0.527396744263735, 0.140662369330878, 
    -0.213569914400005, 0.0186870647370132, 0.574028118982545, 
    0.186966021019077, -0.0487289932596755, 0.0804151894058398, 
    0.368936219983515, 0.134128362329451, 0.0262657914296733, 
    -0.062919798304283, -0.0615117076532272, 0.148240818632544, 
    0.301400543496923, 0.227666320134544, 0.0331242668331541, 
    -0.0537143264164629, -0.159064881051467, 0.317176327246701, 
    0.221030832129489, 0.157800126293605, 0.129456261629535, 
    -0.180646954239207, 0.134636323243927, 0.404136833496106, 
    0.0855372679831303, 0.116187033369439, 0.288837799817939, 
    -0.252387497300384, 0.33289779832566, 0.429337691283175, 0.1737808311872, 
    0.038341861227614, 0.392291701328895, 0.21106193035188, 
    -0.0902754214782791, 0.613492027008483, 0.407744854500401, 
    0.0843281152268159, -0.0251304919663165, 0.13942244013807, 
    0.250289626812875, -0.100274344421366, -0.112829742302937, 
    0.0387531288216813, 0.157275370794275, -0.0499695794096967, 
    -0.0819333396687762, 0.0361006825074789, -0.00333735636661207, 
    0.0537877401910837, -0.0891099489407224, 0.0397648220970361, 
    -0.068826090878886, -0.0129194591607614, 0.00560581237403982, 
    0.0330316584333725, -0.0558276362571639, -0.0493924908830214, 
    0.353176054844834, 0.19637259764679, 0.0547090828146163, 
    -0.0658687992088786, 0.398175019378349, 0.2832759496597, 
    0.170227518981493, 0.151460622243021, 0.220706157741196, 
    0.0296683728911885, -0.0435108157918431, 0.491046134698861, 
    -0.383524156282301, 0.899637067320069, 0.938571115150946, 
    0.18319911853998, -0.649697481019527, 0.775783972881084, 
    0.525399262029259, -0.153216313535261, -0.150321741641852, 
    -0.179501849049146, 0.0865101864706462, 0.264724214978582, 
    0.145744782987855, 0.30507054479621, 0.376956612901737, 
    -0.0835754217452586, -0.0839851186267511, -0.133020463419843, 
    0.01790408116336, 0.00727528792676593, -0.129424436203583, 
    -0.136708719909946, -0.0572139622360732, -0.00504743020253007, 
    -0.121598828072421, -0.112652327897782, 0.0720606539017215, 
    -0.00557757114280193, -0.0417112171269323, 0.157775309253272, 
    0.139245559151214, 0.104213143705423, 0.156775462066849, 
    0.111744084655072, 0.0342797571400584, -0.0499889635827574, 
    0.0487054503459411, 0.163746037945743, 0.206666483949043, 
    0.21066512888164, 0.14505342417712, 0.0413066034092519, 
    0.132448190683632, 0.350573747412698, 0.099089884054173, 
    -0.0497960088128224, 0.024222483572427, -0.0383658605802682, 
    0.339663455446394, 0.442078160965123, 0.223627211330464, 
    0.40999065742552, 0.418951077037348, -0.219025850378254, 
    0.316620004596036, 0.681581308344356, -0.0461818124770094, 
    -0.0460418209066653, -0.0378822551954124, -0.0435573726531571, 
    -0.0374591342906927, 0.0184180867722355, -0.0354274010074399, 
    -0.0516050182938326, -0.023920850143923, -0.070133533620705, 
    0.0441609775747972, -0.136233147027003, 0.0632862140525845, 
    -0.0740250820006257, 0.0437644515132357, -0.123729271203301, 
    0.0318379203075234, -0.0933376126191011, 0.0173242085003673, 
    -0.192373532130857, -0.0399180893791593, 0.0409891828946003, 
    0.0443560478537175, 0.0508030456967063, 0.080148790848997, 
    0.0604762193697566, 0.066377518434944, 0.167242367901011, 
    0.147148546467026, -0.203341230501688, 0.349706865561474, 
    0.35944154898413, 0.137494039710569, 0.242063486025943, 0.41737290600704, 
    0.153459644982347, 0.0510185310410104, -0.556138890286862, 
    0.237503949778533, 0.922690336838243, 0.124973153983392, 
    -0.352466294208207, 0.0517667641577392, 0.770174180971114, 
    0.208922672099584, 0.0919811015515509, -0.356102074879972, 
    0.196374697310328, 0.391407146727052, 0.627179566227801, 
    0.731220326295911, 0.246187585595213, -0.0446806024257583, 
    0.410568619648068, 0.388460684453201, -0.0838709589516198, 
    -0.27516991707224, -0.128940017540889, 0.438084697663633, 
    -0.0143174957686855, -0.139632065202576, -0.0570817457030828, 
    0.0988809075450229, -0.0313103682079839, -0.119473074623446, 
    0.0470666679492251, -0.0255487486037999, -0.157371385192996, 
    -0.1145833135166, -0.15390820754057, 0.0806158497799997, 
    0.137727060535774, 0.230458282768016, 0.230578510358422, 
    0.0863380484718157, 0.0240673945840888, -0.190538915492783, 
    0.431018281016053, 0.394116765441123, -0.097326642453145, 
    0.638770661895605, 0.348926869955405, -0.00539017019133312, 
    -0.0676744524525008, 0.263982607612183, 0.538475238876007, 
    0.332081641611175, 0.663984978346261, 0.895541218388305, 
    0.202056023567421, 0.126385899979401, -0.232806213561229, 
    -0.067987927352719, 0.211234945501945, 0.953385057265964, 
    0.484108765203366, -0.0917335229814198, 0.747908978978335, 
    0.46104355143526, -0.102169598972994, -0.127482238630501, 
    0.250476739268985, -0.171772967237942, 0.0688715813475198, 
    0.101612990717173, -0.0215510767637434, 0.0418543924835718, 
    -0.14443349956001, 0.154439717515756, 0.0264077773371128, 
    0.0161926882227003, 0.415926253527395, 0.242532554041668, 
    0.102062635697462, -0.216856201100078, 0.175841097405164, 
    0.371419328744175, 0.216618543714245, 0.114797261324004, 
    0.123857828204938, -0.127408741972585, 0.0937088477674553, 
    0.4619291221291, 0.373116054651481, 0.127647340556402, 
    -0.111475873434833, -0.00818328486008185, 0.317046263975026, 
    0.281316440878234, 0.188497233129434, 0.168853407264822, 
    0.235910766314726, 0.196395511506509, 0.156624770389549, 0.169496424029, 
    0.12333850830175, 0.0595835756765153, 0.233306602175207, 
    0.133425702827498, -0.0753683897436314, 0.302846278525417, 
    0.309155402215561, -0.102392236620099, -0.175752506272335, 
    0.376980416486694, 0.540784128097869, 0.275464370422754, 
    -0.0481472521081072, 0.392508157642531, 0.335622961930701, 
    0.0945165154905945, 0.0520623931686754, -0.0417558138538968, 
    -0.103484499935502, 0.247035870067592, 0.155950143188004, 
    0.0461466882506242, 0.246441911724912, 0.216790634469272, 
    0.0421092727976918, -0.036755513368221, 0.0181279844674936, 
    -0.0497726504730549, 0.00890563887670996, -0.0681453968543442, 
    -0.0150158259571031, -0.0227756507579519, -4.85255806349783e-05, 
    0.0516431046640389, -0.0791987027589359, 0.0753077775359501, 
    0.134715525295622, 0.090054609008616, 0.161076404923154, 
    0.0960805778191838, 0.169076808588647, 0.360516789655364, 
    0.21157920916358, 0.0490693983619776, 0.217545306620968,
  0.0358615596330625, -0.127963788809377, -0.0789133907591992, 
    -0.072422524386426, -0.0782922473946572, -0.0853954785914398, 
    -0.0796181774110294, -0.0485483215730831, -0.1318335992492, 
    -0.0268570244772564, 0.315082571558284, 0.037394275859003, 
    -0.164804654252786, 0.302848031907911, 0.363860783904694, 
    0.222940984861439, 0.147999185002326, -0.218610060747606, 
    0.245175306923825, 0.309162650009755, 0.147798024533015, 
    0.31102098675034, 0.411096694487516, 0.0849327700628429, 
    0.0965228782049961, 0.560215892927392, 0.055097691338273, 
    0.351000330928623, 0.974077510210527, 0.177162032697425, 
    -0.0459267353480299, -0.00945975336458398, -0.0238929317769815, 
    -0.0189477913980638, -0.0166900316940607, -0.020461203229335, 
    -0.0119054474043074, -0.0162034033838881, -0.00789566624646007, 
    0.010721045497603, 0.0969051761697119, -0.0422819822372547, 
    0.349553747463328, 0.2589977636096, 0.0791872456883337, 
    -0.203192148570993, 0.118159611667787, 0.442943568690729, 
    0.021298452220258, 0.0487532049367904, 0.188070188076428, 
    -0.311102943140667, 0.316580641617346, 0.302666035260383, 
    0.398459723225063, 0.809029045624525, 0.247289534091785, 
    -0.0661075721981532, -0.127163301058518, -0.320650036755053, 
    0.45270724947479, 0.251681926362032, 3.24991264133018e-05, 
    -0.0407392902656125, 0.014743985989034, 0.0452969848155165, 
    -0.0883837311051558, 0.1514111573842, 0.00932012539801991, 
    0.0145255223827302, -0.0597969836688012, 0.191198513866872, 
    -0.107376112673751, 0.104281954906889, -0.366441992988129, 
    -0.0674427046060163, -0.112860974729137, -0.201797699461348, 
    0.0734841867045612, -0.228027547100622, -0.0232900782736144, 
    0.00632102577514979, 0.0425416465484594, 0.0947906126598177, 
    0.062521250028768, 0.0168915660614602, 0.0804318547487819, 
    0.154942693204051, 0.160576941198669, -0.00836604486817359, 
    0.654993938236476, 0.277010516363214, 0.149686462769338, 
    -0.354575887658699, -0.047168868045877, 0.588827234601234, 
    0.390267974416753, 0.115704974716923, -0.0992384638839596, 
    -0.0457679162061506, 0.428048141376006, 0.203556007297933, 
    0.01019393650854, 0.0614673278298215, 0.354164880188657, 
    0.0861272818277091, -0.0221548734023435, 0.122685241441673, 
    0.177263053556956, 0.0141760905818104, -0.0523566833460543, 
    0.00705398209105023, -0.0827187674494253, -0.0102969962962429, 
    -0.0723803880942062, -0.0423182600481722, -0.04209255317955, 
    -0.0379701957328434, -0.0422660426657003, -0.000681025515585632, 
    0.00720710888821249, 0.0310818118378562, 0.285433670058925, 
    0.133840928317169, 0.027733806042562, -0.122025184843263, 
    0.16978427867164, 0.424457926015054, -0.0605931974814082, 
    -0.0314741305575775, -0.562572753425752, 0.374105985807186, 
    0.671564420822949, 0.251502983880496, -0.388604066748203, 
    0.442457440028721, 0.524703291593248, -0.0776228799237354, 
    0.392220761505648, 0.826754721628482, 0.245028085429416, 
    0.103654087080024, 0.0605420373765411, 0.0687412917629464, 
    0.0963716254194894, 0.0653734069971609, 0.0851490096318997, 
    0.132128010194796, 0.121478698708096, 0.0271452277351046, 
    0.0864191632310299, 0.2467415730085, 0.173629982651214, 
    -0.0307511806396218, 0.228755653820839, 0.421848331591169, 
    0.150438036694708, 0.0880232628844155, -0.212979327765508, 
    0.599363547403459, 0.23777481635394, -0.128053202198881, 
    -0.0445068220669182, 0.729962880075648, 0.234382848571429, 
    0.0925941490235773, 0.259082585721163, 0.0840460182488904, 
    -0.07395993293384, 0.939443568232168, 0.294512442310443, 
    0.0315655609366223, 0.345821136605481, 0.336865316696658, 
    -0.12594032788852, 0.319448896994574, 0.272952674723525, 
    0.195587341035376, 0.392878039748023, -0.0666524473574502, 
    -0.319509803941708, -0.123850500003189, -0.222599921111824, 
    -0.206089733106908, -0.232835780433764, -0.264373609499774, 
    -0.0655537124335716, -0.271543686319023, -0.0119831240185539, 
    -0.25465019234123, 0.0742573201470676, -0.0514346558536046, 
    0.0365707016610824, -0.0411588575742757, 0.0179365826179618, 
    -0.00509537666350871, 0.0892646514280617, -0.0450502857534795, 
    0.110753757119192, -0.00828347603702744, 0.199118421931722, 
    0.0100860677416689, 0.0697766148782762, 0.287100676908433, 
    0.278653751276473, 0.149568173608405, -0.091917125569256, 
    0.408560630478873, 0.184949740317149, -0.384808165055841, 
    -0.0653256943560644, 0.706215151210029, 0.347581846081162, 
    0.256070653252159, -0.410224261423069, 0.631137871791285, 
    0.437734156115757, -0.149002850047111, 0.181502402079162, 
    0.883756618088892, 0.243795370961465, 0.136411576160039, 
    0.477052328914884, 0.106596279525845, 0.0524748238132124, 
    -0.236731450699097, 0.18469345340931, 0.290508525792671, 
    0.309487776792895, 0.269459899235401, -0.02704116481902, 
    -0.167498263096095, 0.0117772568277164, -0.146758573286841, 
    0.0724912240159672, -0.0486126430271622, -0.0489874533251947, 
    0.203057533128178, -0.0234110565867614, 0.00315470861625165, 
    -0.12685030315691, 0.112710201458281, -0.0921731549537865, 
    0.055750194355987, -0.0128953614052695, 0.109459271962382, 
    -0.139413397007847, 0.0781971050507162, -0.209618538226102, 
    -0.0520270955690248, -0.0383791683491497, -0.0083932653358233, 
    0.0276356134217336, -0.0543282048891215, 0.0624781826232882, 
    -0.0138009234940884, 0.00830409514057341, 0.0199056267052969, 
    0.025731610422137, -0.0531215503120822, 0.0601121120507977, 
    0.0909236168316208, 0.100993189124476, 0.166367773478139, 
    0.184716577133991, 0.137323576851045, 0.137935719136179, 
    0.208194411731684, 0.200620550487942, 0.170790880050875, 
    0.241546953980088, 0.242688571530065, 0.178128507618326, 
    0.180676000259333, 0.30812153760471, 0.309179510330591, 
    0.175560963255187, 0.0536492198037026, 0.0708554029576142, 
    0.370172116343791, 0.392662278248647, 0.285876920259214, 
    0.182360473357168, 0.0193014119263016, -0.0913058617974089, 
    0.834935089285174, -0.00326974884487366, -0.249212261556488, 
    0.439314973943288, 0.155879465125218, -0.350748088392906, 
    -0.222618490768553, 0.0528486374776728, 0.0136580227489689, 
    0.15915627055289, -0.00745698097269955, 0.0270535132325707, 
    -0.0873496857511422, 0.0998253072950091, -0.0581537741838513, 
    -0.104890185473581, 0.0706286047710719, -0.15112206849413, 
    0.063148375972707, -0.505821682325825, -0.0860220090940613, 
    -0.179394402481744, -0.18500610208939, -0.188260389086587, 
    -0.0685677899241992, -0.10292121430208, -0.0635780135456725, 
    0.0725923413784947, 0.0545299345100216, -0.032842571398727, 
    0.0729672914614205, 0.182561613504095, -0.0429170355521986, 
    -0.0254236620389021, 0.193753065546051, 0.443141113039048, 
    0.249227037212037, -0.338124057097126, -0.0199137194135719, 
    0.546872971081351, 0.629701268269732, 0.371295820926551, 
    0.158057748724462, -0.421694569589695, 0.369787182395533, 
    0.40048006504699, -0.0326260075802, -0.13683392846634, -0.1018139914643, 
    -0.127128517505826, -0.0266819506905041, -0.216657841201525, 
    -0.156507781540417, 0.0452182555677434, -0.0897926618752046, 
    0.0774001464274557, 0.0133405635797614, 0.125471250568814, 
    -0.059485747258993, 0.079063422086342, -0.0819672722632654, 
    0.0328128195682584, -0.0202729686753497, 0.0651072764486516, 
    -0.100028296288177, 0.0705161417004577, -0.152989998324099, 
    0.0220925277204907, -0.116544304831619, 0.0415652225883982, 
    -0.204028656367469, -0.00692612346246713, -0.0436303217892511, 
    0.057337213003642, -0.191324531685491,
  0.0466434584071605, 0.0560800081088396, -0.0943572274489754, 
    0.0017080027885784, 0.0516691289963898, -0.0020016652034481, 
    0.100343990267544, 0.0431101118065875, 0.086499312420549, 
    -0.0216969632290351, 0.0520716615806409, 0.0783131053999315, 
    0.0982777126834341, 0.147470985083716, 0.169031301683326, 
    0.14156033234743, 0.141317673533012, 0.189313737124555, 0.18145063905056, 
    0.176363908440371, 0.192703256376165, 0.058708262199859, 
    0.133921334657042, 0.506265707983929, 0.230310942791856, 
    -0.0400997918768876, 0.0642336003678176, 0.539508414976373, 
    0.226022267791872, 0.0716647686037721, -0.0887191965395647, 
    0.0583708934762593, 0.124826123469575, 0.476019523550144, 
    0.574301505403067, 0.110763183723172, -0.30532327723008, 
    0.10666840838143, 0.568848043579342, 0.109375209880943, 
    -0.0671020809967359, -0.0369388575930469, 0.0690195519302978, 
    0.389909776955701, 0.161179760394062, -0.0696048800296294, 
    0.228653532391098, 0.222710636769555, -0.107296581626392, 
    -0.0543325081823902, -0.0931065398797638, -0.253860033105957, 
    0.134521874337485, -0.061287744865144, 0.0971160604663423, 
    -0.226466498895831, 0.0359714359306045, -0.171322552071667, 
    0.0319249497564491, -0.262480208565864, -0.0173738225459496, 
    0.0238254295455498, 0.108262991200534, 0.166187459399191, 
    0.117048077332143, 0.0265336823791278, 0.186632530382126, 
    0.297471881005005, 0.0271135409556767, 0.00312604835845329, 
    -0.25297240955514, 0.449876339915169, 0.408084962124564, 
    0.0862824221213554, -0.199570737616339, -0.106382879994496, 
    0.548633260432038, 0.422284068908665, 0.134546161076018, 
    -0.313777597360603, -0.121370399100699, 0.507637616151206, 
    0.644966236915571, 0.174573281724581, -0.267020101107982, 
    -0.0892552530049911, 0.479112015044817, 0.542978307554058, 
    0.314272094815272, 0.408191047985473, 0.612324179517715, 
    -0.0127332909570982, -0.0697746987705559, -0.0244657822798662, 
    0.239708343742924, -0.301911893520982, 0.115477096284859, 
    0.240597641752003, 0.40398990332677, 0.381788104512328, 
    -0.0135894377182104, -0.0831311321977299, 0.126046689634355, 
    -0.013552936409337, -0.111650501600583, -0.0160154768654001, 
    -0.132994756367937, -0.0904615286265559, -0.0261025254866962, 
    0.00444104134134708, 0.191086360044677, 0.116727232747364, 
    -0.0265669300078194, 0.270932028015389, 0.191024763874055, 
    -0.0284058889986274, 0.203673820323537, 0.345045413103821, 
    -0.0071927192022322, 0.188965133309913, -0.208596601517866, 
    0.503958469650063, 0.319991133172183, 0.30563577424884, 
    0.399160097062626, -0.3112591287245, 0.553759943478239, 
    0.608562345541333, 0.0457831564131265, 0.548963557621976, 
    0.77557902131659, 0.00867891412038939, -0.296542293721435, 
    0.234194148189151, 0.418367666965011, 0.0314866261197316, 
    -0.184937721072982, 0.5154078225765, 0.507712581263552, 
    0.304413625030456, 0.300487541208226, 0.269677376947672, 
    0.121136231710772, 0.0761298026782096, 0.0845980416305218, 
    0.0398650627012573, 0.163051031926352, 0.197391488578781, 
    0.0603142465889393, -0.0254898942664151, 0.291840006208856, 
    0.25643510921876, -0.185440861524731, 0.437193017141568, 
    0.38696120318787, 0.0639434273323351, -0.200260363947926, 
    -0.0439208961219078, 0.491195566807394, 0.297378046857289, 
    0.067437789628954, -0.0451660752213511, 0.0704864240886204, 
    0.442544837786156, 0.0642788534024265, -0.0971107418215486, 
    0.00340133623978872, 0.362653233311305, 0.0882631442919939, 
    0.00364786964492275, -0.194379893928332, -0.0442966146110377, 
    -0.153335783240549, -0.113568947599838, -0.0532497259560241, 
    -0.135354034566307, 0.0116523689279978, -0.120771136215934, 
    0.0366167788175857, -0.13922891804097, 0.0192244460408457, 
    0.0407764600074611, 0.126028960263616, 0.169245700561101, 
    0.10100536099084, 0.0283677551920487, 0.140617479314275, 
    0.379260041947344, 0.129945504452801, -0.275524750987524, 
    0.0666493212749924, 0.552349334854405, 0.188133130191222, 
    0.0636961461095119, 0.120815469500807, -0.0965112947904398, 
    -0.143513798568825, 0.707638540990478, 0.435366141392131, 
    0.107121414805816, -0.00582225069488097, 0.17282013257613, 
    -0.344029931388823, 0.44310308408793, 0.386958474098366, 
    0.044795207461567, -0.28915755433537, 0.185022981784565, 
    0.265558018605891, -0.0283098964812715, -0.0675427916208849, 
    -0.287219823888723, 0.0734438269233366, -0.0704650122133153, 
    0.072322059543003, -0.154383651001707, 0.0479796899015629, 
    -0.0930509739065914, 0.0366464104075036, -0.302868246070403, 
    -0.0343290745161514, 0.0785850924545294, 0.0929351892445472, 
    0.122503048152804, 0.165877701817225, 0.166293583698089, 
    0.20013104552499, 0.221955864287721, 0.127752842632476, 
    -0.135509707454945, 0.419955673652461, 0.393311632758861, 
    0.176052188895622, 0.189052046199704, 0.155452392738581, 
    -0.0360044013981462, 0.744330874564164, 0.485132165089711, 
    0.083522346376888, 0.145897324391656, -0.15715766608315, 
    0.667842528251192, 0.0146389806667513, -0.0887219842965248, 
    0.138445999716755, -0.192522889612764, 0.786627483023973, 
    0.268134703354823, -0.06396965011866, -0.0643864413111168, 
    -0.181909415874332, -0.29559242340472, 0.0334469108137981, 
    -0.315235602340771, 0.0361134571648079, -0.316945285962774, 
    -0.00394835694125058, -0.283431529941957, -0.038071196832209, 
    -0.200535414177767, -0.00321831736945331, 0.076610721447868, 
    0.126842994033222, 0.146839099764163, 0.145539331645846, 
    0.162068661810276, 0.183393878651497, 0.165684086324794, 
    0.109500587594575, 0.0976571724033594, 0.130430201898454, 
    0.139946969312673, 0.146655758103088, 0.193834291108625, 
    0.221858075399218, 0.159217128801618, 0.134024317181978, 
    0.29369818003889, 0.209985592173365, -0.0569335016564692, 
    0.428002815178949, 0.349725436267888, 0.0533158435945193, 
    -0.213010403724029, 0.185108094718777, 0.553846225650357, 
    0.145479276880481, -0.0305600657908538, -0.0419130502251456, 
    -0.122613728753499, 0.267088465782059, 0.642753607429823, 
    0.152507930354824, -0.208105158981124, 0.246692191064424, 
    0.302529874019554, 0.0036188258229596, 0.143939279508965, 
    0.724300484006747, -0.127896125181135, -0.128642329251609, 
    -0.0207903185037782, -0.0917378242496148, 0.00788227006009352, 
    -0.202778827560536, -0.0472982351095797, -0.191643338204923, 
    -0.170103889192386, 0.090988377022543, -0.212635270569272, 
    -0.011173014300379, 0.107757191801433, 0.194186409189664, 
    0.217399265227011, 0.185731322560501, 0.171579940384227, 
    0.294384348725583, 0.414150831944643, 0.318977559645099, 
    0.165772573115005, 0.142158454465021, 0.391328340254255, 
    0.466374842523941, 0.287099369532697, 0.319599013876385, 
    0.632637081741027, 0.482252504391096, 0.17267622839753, 
    -0.0700000995364356, 0.478847835394992, 0.593108141127753, 
    0.130387335075425, -0.0872915539082742, -0.0619957988423457, 
    0.365128670359922, 0.509533844881408, 0.246614346686141, 
    0.0318222325221394, 0.35380551425509, 0.243077782442869, 
    -0.0440923786020395, 0.206523821447115, 0.107833576176511, 
    0.647380444169107, 0.8066690396122, 0.090542144904114, 
    -0.202410130686506, 0.414026195806442, -0.114244853183975, 
    -0.211811213796992, -0.333537742552385, 0.159162488613178, 
    -0.256748935577124, 0.0477808532890324, -0.266444283683315, 
    0.022367190678625, -0.257134392385682, -0.0186966465166822, 
    -0.256841163740235, -0.153907419752214,
  0.0566637824666357, -0.0353456767880599, 0.0983568416977215, 
    -0.0870092100648161, 0.0590355260851567, -0.201227846544766, 
    -0.0353625889236151, -0.0935883139655669, -0.0928323209059453, 
    -0.0478089375458732, -0.0110519490260741, 0.0565593079525605, 
    0.0183211791306472, 0.0377952847950131, 0.0341801150139238, 
    0.0360350222493415, -0.0234224742848493, 0.0255917386032968, 
    0.0266484505995883, -0.0204889353743734, 0.096712452196632, 
    0.0720821454219601, 0.0883136302712993, 0.290686512755497, 
    0.17565365671748, -0.0474537283960953, 0.29662656814791, 
    0.288887324334273, -0.110791749981134, 0.141871822985682, 
    -0.0549953923300773, 0.703027823461687, -0.0466771507142259, 
    0.00226593712499987, -0.426324968040982, 0.419097998685957, 
    0.582107143709291, 0.342599720096481, 0.314285581659703, 
    0.260429896165556, 0.066420641908643, 0.323584262132644, 
    0.281235501702162, -0.0133348318535991, -0.141310273508745, 
    -0.188548058525944, -0.0717666348868972, -0.0285530766293919, 
    0.19711372282534, -0.23905638286257, -0.0233866687241794, 
    -0.283281291257912, -0.0337312745214969, -0.126654828317886, 
    -0.0045141061386294, -0.0742955036839586, 0.0328440480523054, 
    -0.134097886520551, 0.0129753947076847, -0.435686525910511, 
    -0.0621545833216453, -0.0364085156645002, -0.0154955751869555, 
    0.0290376583934719, 0.0117007293036954, -0.0380207864121537, 
    -0.00153887474496814, 0.0537054409863504, 0.0770443400855308, 
    0.231495475955635, -0.244873752733924, 0.353011919886303, 
    0.500496592076969, 0.119799297223764, -0.224497826311586, 
    0.168417723385391, 0.0892176351699272, 0.750160248439073, 
    0.592024552273746, -0.0255293937529214, -0.132439655236456, 
    0.0791248295912555, -0.0749071191304826, 0.0987882854036486, 
    0.0536031281198985, 0.0294813944635286, -0.0263518425043195, 
    0.113080102314663, 0.240725441427557, 0.0151662710376948, 
    -0.102529195913928, 0.0021723302075768, -0.219740236075834, 
    -0.00767106378235895, -0.0907799246420362, 0.0608515679392785, 
    -0.308113763063301, 0.0105258384958136, -0.298161613546604, 
    -0.239626262992997, -0.00765973029730262, 0.0460258394932029, 
    0.0819233488974469, 0.14011128301946, 0.139208658239321, 
    0.0830236935768698, 0.134133378771395, 0.268679277369774, 
    0.157959297878251, 0.00574128289396037, 0.145109058709433, 
    0.349340447104124, 0.222063658609257, 0.16548716455545, 
    0.527224539039128, 0.35322115666808, -0.025451865734456, 
    0.37058548245225, 0.696551674635091, 0.142215878065903, 
    -0.123696871976906, 0.157927001709839, 0.898467992094485, 
    0.0755903941439498, 0.137496089375974, -0.259107535049517, 
    0.103757365253683, 0.63418406858373, 0.349574853892144, 
    0.0821126615279106, 0.0572397631015029, -0.099281512130081, 
    0.623742316162197, 0.226777890380632, -0.0639355624251853, 
    0.174025285097138, 0.201406548527934, 0.393860720838153, 
    0.304353582376307, -0.236288176857918, -0.328548920557541, 
    -0.139864493626792, -0.239074533734191, -0.199537151990438, 
    -0.277712693677703, -0.155495900227296, -0.264120852301474, 
    -0.201103597341196, -0.213105714950397, -0.110768739390449, 
    -0.0906152665119586, 0.0154573596857241, 0.00742032982940084, 
    -0.0226218609050065, 0.0222343766345899, 0.0706007094172852, 
    0.107853705930709, -0.0227072849525757, 0.0560798650713278, 
    0.061540125792682, 0.0615120636041642, -0.0415430091199235, 
    0.0214994313021914, -0.0170263306118572, -0.0260669507601979, 
    0.0615765295345868, -0.0288243560208032, 0.0210409000925205, 
    -0.0241359790770436, -0.0400303363009437, 0.0363180774702138, 
    0.0915504812964802, 0.100317036805605, 0.0935303585119745, 
    0.102907862624745, 0.0983579136133138, 0.105243212442777, 
    0.129079492876079, 0.106907696653181, 0.0634527269905344, 
    0.134240348411565, 0.16497825178064, 0.150714491217318, 
    0.222194412734868, 0.267530307906753, 0.150872536417591, 
    0.127677923505702, 0.390585239839106, 0.204406188775838, 
    -0.078053734402554, 0.28645149336998, 0.410103299327901, 
    0.153671981516404, 0.212448528386945, 0.123051689427203, 
    0.965503642929208, 0.757027133076038, 0.138488793517592, 
    0.0513501021422458, 0.131960871657749, 0.373792855012893, 
    -0.0696122414423951, 0.83155985343715, 0.521800301569997, 
    0.169548438694906, 0.203023687270842, 0.153342442254267, 
    0.591025239271806, 1.17116342012236, 0.0227896645024999, 
    -0.219567912876103, -0.367446355894478, 0.135098864001616, 
    0.0194287407326802, -0.0660031003480936, -0.0631141246271224, 
    -0.0675775665870915, -0.0908043482489883, 0.115534090901126, 
    -0.0347523223013493, 0.0226290999756056, 0.155481436720978, 
    0.144078758131299, 0.0332660780065804, 0.0673658466517338, 
    0.0604620540885404, 0.055158361210626, 0.28501333503614, 
    0.202960646312135, 0.0847581634346105, -0.00650423021353544, 
    0.285056416114858, 0.3075043767577, -0.119855079399142, 
    0.0400975547439066, 0.72037941777723, 0.190525443616732, 
    0.0796595647577037, -0.166126754882906, 0.241486045655089, 
    0.445333260204592, 0.212799764375624, 0.060665959076371, 
    -0.0340250827557235, 0.393044847176162, 0.284875416753883, 
    0.0355707713436185, 0.404714614455145, 0.519701782434647, 
    0.111957572945016, -0.137263078131029, 0.0146522463007798, 
    0.655436086268894, 0.186565715238473, -0.0516336895451518, 
    0.0423790849897654, 0.304020384876015, 0.298960692819933, 
    0.331224488032843, 0.374080483405992, 0.537204397278029, 
    0.327882038954313, -0.200098991359067, -0.429818703946861, 
    -0.311779317546417, 0.29580867435013, 0.458367825606467, 
    0.823440999651172, -0.0744492957125606, -0.403402655361421, 
    -0.510354039537078, 0.135110480210146, -0.375613776633776, 
    -0.130276976967856, -0.200825357404933, -0.185682990299401, 
    -0.197826280316661, -0.163347258951739, -0.195675704984886, 
    -0.0603253692639149, -0.0853140171648777, 0.165247580850982, 
    0.0621009466071411, 0.0992077758082886, -0.0491264857592648, 
    0.0662963075042871, -0.126810377645957, -0.0305941453488217, 
    0.0361074898408291, -0.0612835211724505, 0.228847252234326, 
    0.0220036364670419, -0.104174960282341, 0.390768114154477, 
    0.245185531084489, 0.02435918044137, 0.430406078715386, 
    0.318103607693729, -0.0742710718405668, 0.542486904243072, 
    0.439303488126323, 0.0917738401372169, 0.535827058308304, 
    0.267554795176085, -0.225698140370769, -0.0569198662605817, 
    -0.169157137235158, 0.587326756306616, 0.17789629617248, 
    0.325570593509221, 0.60683030209187, 0.243548203204304, 
    0.081642067459279, 0.0482386203618862, 0.0573208700420512, 
    0.0617310927130987, 0.0650954653240555, 0.104757336863279, 
    0.0479675196224789, -0.00639711390228008, 0.0118585632731173, 
    0.0398680992788421, 0.094627288371494, 0.169291194869852, 
    0.308637859981822, 0.452517595538772, 0.261312953259998, 
    0.0174175371524189, 0.475426016076771, 0.266904991109613, 
    0.166319058681878, -0.264321169951751, 0.471713592235867, 
    0.522043187508985, 0.138945646983639, 0.0473480935429452, 
    -0.249634096554385, 0.500070860525406, 0.332107767111811, 
    0.0187320148181117, 0.483515707423627, 0.501748008929327, 
    0.162902840689588, 0.0681733074610056, -0.0425366919958858, 
    0.223946946657019, -0.0422712058999407, 0.526234512344138, 
    0.284636112714543, -0.169213604472498, -0.154080991185889, 
    -0.0970294976848778, -0.109297711593154, 0.0108526522175194, 
    -0.0581824623097933, -0.0020693658971517, -0.000331086857056226, 
    -0.184326844163481, -0.0076083467314898, -0.122211719641922,
  0.32056355106826, 0.184536061435452, 0.0798514974416896, 
    -0.0861313998156578, 0.225100148776179, 0.319486591752609, 
    0.141044228930399, -0.000135403245685492, 0.297133563336587, 
    0.259480133974588, 0.077217761873471, 0.0472521189045076, 
    0.0840008225476202, 0.0906635210505992, 0.101978895487671, 
    0.068287369319374, 0.0103276699284263, 0.194598592278733, 
    0.139189833362055, -0.0698228253332732, -0.0752251952691879, 
    0.229805216735927, 0.342619506542923, 0.421165428883445, 
    0.182282820733627, -0.191193128348012, 0.0728678480336878, 
    0.549306127797323, 0.0168292546623164, -0.0943153105422896, 
    0.259660833479784, 0.537468944867642, -0.111462393286877, 
    0.480643115294925, 0.559168615884647, 0.163112337374691, 
    0.679949241819426, 0.811216444175603, 0.490100590608917, 
    0.289228538781515, 0.0494650789380461, 0.355180139529477, 
    0.181986704265599, 0.195738263022883, 0.185882190306443, 
    -0.145031025858246, 0.234741492905442, 0.230504813496777, 
    0.0542709961330337, 0.0244496666373877, 0.209233637567385, 
    0.199813576282485, 0.0735799387504613, 0.0172592811004924, 
    0.151411416311252, 0.0490906437009341, -0.10317723455177, 
    -0.0546354557260322, 0.257253901894742, 0.0855687451320175, 
    0.0261610415679405, 0.090489629398026, -0.0186167012221822, 
    -0.0259421587699212, 0.00769386340867806, -0.0244960859696309, 
    0.0450076423593848, -0.020413685237811, -0.0100527718032359, 
    -0.0266396466768052, -0.000542671799690544, -0.121383071760281, 
    0.0330776401646859, -0.0498122170723191, 0.0256415875346102, 
    -0.0889876489092945, 0.0182662648296721, -0.0773904044652313, 
    0.00511327692679657, -0.136330868679765, -0.000384806333295046, 
    0.0339271470198816, 0.0698857116954236, 0.12765325379339, 
    0.210633218172106, 0.154682164887936, -0.0725185952613182, 
    0.365533863658374, 0.0442863286746714, -0.195071526709982, 
    -0.142284980225529, 0.672585520831843, 0.15305924217325, 
    0.0314273915947487, -0.0969641387686831, -0.186557878443981, 
    0.375602579021574, 0.689764635212744, 0.217756076634191, 
    -0.0648745384082615, 0.257257852340851, 0.374707402111455, 
    -0.261763960367422, -0.0897755938547689, 0.0235439961222103, 
    -0.127642374699709, 0.233259751287113, 0.615155922258206, 
    -0.0223945210620841, -0.108731955913046, -0.199908282016425, 
    -0.193781883602512, -0.0820203603985138, -0.285733964752953, 
    -0.10334561806309, -0.201326614749224, -0.206988420487279, 
    -0.225959080097434, -0.131840696690191, -0.232342722944798, 
    -0.0600619359499707, -0.103799117257374, 0.0805968817041214, 
    -0.17307176075958, 0.123850718753331, -0.0494645953540755, 
    0.0338700110565942, 0.00979167988334231, 0.0596208653712293, 
    -0.114707301633349, 0.0309845375637401, 0.0555569024850388, 
    0.0612190461426364, 0.0498652867317967, 0.054743680906186, 
    0.0426359814201538, 0.0487199594743129, 0.0728294771364991, 
    0.0559994357303111, 0.00932217029358347, 0.0715713917880826, 
    0.115307036978193, 0.155782737722402, 0.158820477075788, 
    0.11866176918146, 0.142660401616177, 0.249912078801775, 
    0.219472792017866, 0.134951868227645, -0.170200919830029, 
    0.425783127599874, 0.295676828044655, 0.00315281977598064, 
    0.297396509037289, 0.381427720425815, 0.06008745223938, 0.50121539073182, 
    0.593076890244572, 0.147856833483401, -0.120621617342924, 
    0.633009616146472, 0.324602813692435, 0.0436647251161157, 
    -0.0462342768445881, -0.246789742945725, -0.325774886797974, 
    0.214325575508513, 0.405347160664976, 0.434801260128991, 
    0.138489709822448, -0.278379335787117, -0.243588396006456, 
    -0.242786225225801, -0.0623329026739487, -0.23922707201072, 
    0.0300481910605833, -0.242093627708884, 0.0408203786332721, 
    -0.321367595855674, -0.123013602880404, -0.0112384664136182, 
    0.102046282163944, 0.0389509130082378, 0.0789209731077823, 
    -0.0269103227040832, 0.0140235750746731, 0.0590634876794707, 
    0.0311992590455501, 0.0933213374489174, 0.00346398192902245, 
    0.0491751420337767, 0.0919325554531688, 0.122206196297694, 
    0.153844268798292, 0.184331155537238, 0.175658105910022, 
    0.137409160187722, 0.13522032239314, 0.205286735409327, 
    0.219708871750097, 0.165640725987625, 0.136350538183433, 
    0.135129318560183, 0.128431378574803, 0.125002686409466, 
    0.121915652684116, 0.134231195098317, 0.188790425935379, 
    0.171186242614254, 0.0717903670128314, -0.0538280702326611, 
    0.241470093095937, 0.369180208245987, 0.153149138636651, 
    -0.0435755449246759, 0.294843122315846, 0.337296811992439, 
    0.179784829728119, 0.275315353881103, 0.311154180957416, 
    0.00132733678287892, 0.799209768946637, 0.56149148986417, 
    0.315365361276336, 0.209116570660451, -0.375790608889892, 
    -0.0176352233552691, 0.593470035014446, 0.490848923883082, 
    0.264680421608206, 0.0989512593763787, 0.389600862543592, 
    0.0273652551962753, -0.0488375321027727, 0.0178024770752265, 
    0.110441875411453, -0.121669301118283, 0.095485106117583, 
    -0.412037707334456, -0.135715526944568, -0.321483818081939, 
    -0.122401331100187, -0.276480006668225, -0.200843364544511, 
    -0.0819283786715853, -0.236992674004747, 0.08435718580931, 
    -0.183995974822757, 0.0946711903954797, -0.273857406552142, 
    -0.0342565065168211, 0.0187856322219171, 0.0530461046246848, 
    0.0875739753707274, 0.0653411977931894, 0.00276288176856161, 
    0.0611281325245096, 0.219646548783363, -0.107924316606227, 
    -0.221079315950287, -0.0538535704906435, 0.50814564457304, 
    0.0948363794847551, 0.213040984641522, -0.553018637522818, 
    0.32370749808107, 0.596162675848425, 0.205712041898489, 
    -0.0300973928891937, 0.427968068524542, 0.231721387496479, 
    -0.231670896420871, 0.135233391287435, 0.610854922017247, 
    0.0693394398569365, -0.0516641422463682, 0.227791868648937, 
    0.139070297543498, -0.0918791130678698, -0.109844067822077, 
    -0.26631108365347, -0.25827992088324, -0.0166486569949554, 
    -0.0513482144870652, 0.100018709142136, -0.166566730055305, 
    0.15203267388654, -0.0968444246855514, 0.20218037201578, 
    -0.0944819204271287, 0.336995450752851, 0.142633165688012, 
    0.645353703749809, 0.288625447368771, -0.0882428622066474, 
    0.138569793248312, 0.617186057206912, 0.0335277869834852, 
    -0.0115039296056445, -0.138628411422337, 0.0641736134732992, 
    0.398850717957423, 0.396656320322538, 0.309735261774797, 
    0.328227688553016, 0.326010903561467, 0.200487637348984, 
    0.15274278446452, 0.358026779455008, 0.278433276327076, 
    0.047128919211782, 0.0182260739466203, 0.0339498649649406, 
    0.0309964524347856, 0.0341516597206276, 0.043772774696608, 
    0.00845085095420456, 0.0557278371022875, 0.0673703295312188, 
    0.0215609926437191, 0.234759640833039, 0.183491796085235, 
    -0.188474210280551, 0.321755644992551, 0.416422838370345, 
    0.197538295090522, 0.0997612475142527, 0.0400324350363459, 
    0.24632341852206, 0.439081698171344, -0.0019092031349606, 
    1.30482787567334, 0.0499446573951973, -0.453932055777597, 
    0.0391466174103788, 0.733574208070221, 0.319042641306917, 
    1.0692595404383, 0.659095641855644, -0.0640706076750086, 
    -0.0991407401116058, -0.0656873602064711, -0.0731742396851492, 
    -0.0342087112589988, 0.027756163281074, 0.0568655328663973, 
    0.00130425998797558, 0.0273264517285457, 0.132194319871486, 
    -0.185233992609575, 0.148341546073691, 0.257829269264436, 
    0.101883857261269, -0.0226764948809867, 0.0940953204328292, 
    0.272391148653905, 0.289777159212193, 0.121736074733112, 
    -0.0855529101969251, 0.0402647969792598,
  0.220246858653555, -0.0852522067261885, 0.223493201247918, 
    0.39018475986737, 0.124330561540249, 0.0284027832005635, 
    -0.184826606303182, -0.0820275474561215, 0.354879569271581, 
    0.466641549817052, 0.352581866306116, 0.201599465586157, 
    -0.110065632540211, 0.738974821148582, 0.255186831883357, 
    0.14632662708506, -0.405603314863304, 0.747846706715574, 
    0.444200876049424, 0.0500457318121143, -0.102549190200574, 
    -0.289405208472797, 0.307410194767525, 0.671399387501017, 
    0.236937588850658, -0.0281972786697476, 0.309645916238203, 
    0.296766157537551, -0.130757213191956, 0.463617748918087, 
    0.724797369074735, 0.314931339648471, 0.115251267874495, 
    0.0187591435668431, 0.447135321596403, 0.408998474757319, 
    0.0552534419914476, 0.289551740246267, 0.716151423191613, 
    -0.0851721483377938, -0.0908049616834332, -0.0447092880695765, 
    -0.0397821357678098, -0.0528559071800866, 0.012808963147146, 
    0.0138150694717445, -0.0247159721340518, -0.0396596357243345, 
    -0.0127728411804148, -0.0409311052795914, 0.081457090188988, 
    0.116765883999105, 0.122759305384483, 0.127742521088849, 
    0.117855462603249, 0.103807488849309, 0.133301388453372, 
    0.156063618936508, 0.183385020991421, 0.128924753467672, 
    -0.182089918572898, 0.0349601518145639, 0.470660024148919, 
    0.258033590113727, 0.0823939441310242, 0.189595411754859, 
    0.371379348023363, 0.138385962980194, 0.466633262457154, 
    0.682398207378091, -0.0409270385333172, -0.0896450279920479, 
    -0.582020493701855, 0.147940208626899, 0.951843719791932, 
    0.214318574405469, -0.0748089776713005, 0.527561324389292, 
    -0.290862554078826, -0.402417865449283, -0.232795035538241, 
    -0.162340396293643, -0.21930114625039, -0.239850737245709, 
    -0.192424175087248, -0.146979443258352, -0.251647476439614, 
    -0.118601654383425, -0.164445195172354, -0.17155756473856, 
    0.0241334904775237, 0.0736040289923336, 0.0743270837071507, 
    0.0669965338633869, 0.0915658065532121, 0.0677878889010199, 
    0.0962208463200873, 0.0967092143509988, 0.114084254483425, 
    0.0681601406320936, 0.0966196694507847, 0.114884247607482, 
    0.120920236582916, 0.142357411348936, 0.16126129688201, 
    0.143213246953427, 0.146896331540321, 0.130856404910259, 
    -0.00393071093743878, 0.18459543133771, 0.398603647007975, 
    0.116607056933297, -0.136277647410711, 0.123059013259457, 
    0.374675667825296, 0.351860722254347, 0.355070908785872, 
    0.325087232126419, 0.207067267651493, -0.301223859537585, 
    0.532926504430375, 0.334792027468354, -0.166444527712309, 
    0.323965575295539, 0.73607736621053, -0.0471163141844115, 
    -0.34628413910708, 0.115815024339638, 0.38078450928818, 
    -0.0205891274562777, -0.233195376036384, 0.175089705526934, 
    -0.171353647613494, 0.14545157825575, -0.242902368261162, 
    0.0890805148823396, -0.218463520038956, 0.0119449328651391, 
    -0.316870204604758, -0.150026260851027, 0.00705663425549718, 
    0.104627502550209, 0.107822993174753, 0.121266467739122, 
    0.191373007610192, 0.174848903298994, 0.10281183919593, 
    0.138527341512348, 0.098320314813031, 0.105732136391318, 
    0.0452219833067656, 0.0554334820909921, 0.049766790526683, 
    0.0471512685570545, 0.0958258926445441, 0.048298491840881, 
    0.0614190127381768, 0.0804263554618363, 0.0768515061874031, 
    0.0214050512559127, 0.0643062504978252, 0.0930165002186114, 
    0.112697906143776, 0.140642377705957, 0.143980911388473, 
    0.116013823211707, 0.141776655842154, 0.216474518164908, 
    0.133158668296547, -0.050552438434986, 0.212979560517526, 
    0.38610383792837, 0.144743901585004, -0.125211862622215, 
    0.175098508398622, 0.434501104442602, 0.300520943278995, 
    0.187674676955543, -0.0359053064085343, 0.559028851009593, 
    0.179960125660248, 0.0539443970912064, -0.24631122752559, 
    0.299243395303448, 0.422149736610091, 0.270312864315717, 
    0.355066505552334, 0.381660927828962, -0.01049190759301, 
    0.422151615395849, 0.29232302479217, -0.12312650939816, 
    -0.112814455578402, -0.0639223642526478, -0.131230910434045, 
    -0.0353471353688597, -0.0270843051986784, -0.0136050541606839, 
    -0.0557496905714653, -0.134775153640738, -0.123549580214929, 
    0.0845751957904904, -0.323201690037388, -0.0635489123959368, 
    -0.177221009508582, -0.27901246164046, 0.0645327443276128, 
    -0.0910049701547234, 0.0099585914618725, -0.274942549611851, 
    -0.0506224988962561, 0.0235417574169461, 0.0770016206164682, 
    0.130157361066284, 0.0892071357198184, -0.0334996054117133, 
    0.0468207364860506, 0.386879404043582, 0.036922286053376, 
    -0.321385985351304, -0.173196848910657, 0.72628068034373, 
    0.300567743068709, -0.138446815808754, 0.151974726552698, 
    0.624819766831919, 0.604295061036511, 0.293191275725505, 
    -0.0351990582580076, 0.608889964185547, 0.188880962292403, 
    -0.266327975533865, 0.000436333546069742, 0.809806183119798, 
    0.0737950847663947, -0.0786089890125074, -0.090925897394874, 
    0.481969392366521, 0.376298346506141, 0.148956546472748, 
    -0.0184589923709377, 0.209077672988472, -0.0118057645867412, 
    -0.048456620613679, 0.0260961477679776, -0.0512618236931347, 
    -0.184208300603633, -0.292721037293078, 0.0220930707771764, 
    -0.0298856331236842, -0.141552130027993, -0.0367569178750457, 
    -0.120787267037891, -0.078292591209264, -0.0708097400710776, 
    -0.117396132272697, -0.0308719000030206, -0.105612521648614, 
    0.0198655560922592, -0.0924864882807959, 0.0488619817515286, 
    -0.00842180560298884, 0.0362509612959802, 0.00897530745356698, 
    0.0337555790058957, -0.0133809525623043, 0.029910785847163, 
    -0.00323324701046981, 0.027929239908519, -0.0256019191514291, 
    -0.0396434797321502, 0.188406711724521, 0.17387969671987, 
    0.0852836208689459, 0.109079254976637, 0.0705663915474963, 
    0.339868763936699, 0.297629780429267, 0.0135151593909413, 
    -0.049564454510951, 0.474084003027235, 0.474181979493653, 
    0.469839154958805, 0.114279405326098, 0.366523049775686, 
    1.22891399764431, 0.183309089249882, -0.0397225099531182, 
    0.0999260661544475, -0.112999125915558, 0.00486725827279036, 
    0.307358675775673, 0.0797168857005624, -0.00630638404405343, 
    -0.147216062232333, 0.106552099735037, 0.0735603576140063, 
    -0.0268347773146804, -0.132095314628447, -0.0504000223696939, 
    -0.189552924218565, 0.0918079951806709, -0.207012872761522, 
    0.00374350098318371, -0.144910325360942, 0.013532494978068, 
    -0.118155904329078, 0.0498413205767262, -0.161194548566194, 
    -0.0202622394281386, -0.0187665032468436, 0.0160734297599157, 
    0.00367053376768824, -0.0360308512514323, 0.0414735915485385, 
    0.0202833504365061, 0.0418502627246136, 0.0516619963919037, 
    0.0550679986094955, -0.0267068268017789, 0.0771673190858027, 
    0.106737732606557, 0.0907669346930562, 0.19049324315676, 
    0.19754426076835, 0.0492264746069933, 0.186858012723881, 
    0.363996597804382, 0.0331263395737739, 0.0883259440439506, 
    -0.166220780408552, 0.454741564042627, 0.262431452743985, 
    0.0119193457701814, -0.210440069796537, 0.304504070933831, 
    0.847556420657563, 0.210929552727675, -0.122609027281403, 
    0.154643753322315, 0.482407794463941, 0.107206088549467, 
    -0.112644873807416, 0.297288960954232, 0.264952769736003, 
    -0.248747475812973, -0.391542834877932, 0.173610275977092, 
    0.136684920943384, -0.177194894487841, -0.185949094636777, 
    0.0789737218753864, -0.136128325646631, 0.0347590764637593, 
    -0.227835870865914, -0.049894705377192, -0.106545441646708, 
    -0.141123133052949, 0.0826804003336175, -0.131524164351092,
  0.242671282917082, 0.218372525199344, 0.188625654045269, 0.190329571466969, 
    0.199234471912244, 0.202612465565621, 0.234121965718834, 
    0.199551053795911, 0.0876302672383775, 0.158605009269837, 
    0.410537390381908, 0.213265719938634, 0.000673468277153519, 
    0.413120206247342, 0.381975106011713, 0.1676048774287, 0.18016313257759, 
    0.0696595428528248, 0.23887748834515, 0.786411075642182, 
    0.237033967436285, -0.0571440888728535, -0.3215565837535, 
    -0.149099108444927, 0.603359988215013, 0.377732100165705, 
    0.259687952314815, 0.280849996059742, 0.152853626897378, 
    0.544664665173323, -0.128024136917347, -0.110913535423648, 
    -0.123545547135092, -0.125814167625811, -0.0894488440574397, 
    -0.122485978785715, -0.145006700499176, -0.00654633692474638, 
    -0.160732377550524, -0.104900215251089, 0.000256338473923437, 
    0.0450168666608545, -0.0798800020588033, 0.000904069236504379, 
    0.0317137978365767, -0.0425285938094093, 0.0189592500683819, 
    0.0765679641168704, 0.074424411564304, -0.0370398683842401, 
    -0.0675061367618032, 0.120617933970318, 0.214744909057602, 
    0.212636363658833, 0.322791035759198, 0.137465937773952, 
    -0.142870535180337, -0.0527834240645601, 0.298410876274599, 
    0.266268242201954, 0.385958617497691, 0.193069667773613, 
    -0.342348761876915, 0.33741212559425, 0.170019345279748, 
    -0.257473187612602, -0.645310556062255, 0.225961255025845, 
    0.198887411753083, -0.30772049670925, -0.135340676230089, 
    -0.0320452411664489, -0.131612940614629, -0.0804444138991182, 
    -0.10587932814653, -0.0720734589402737, -0.0976460331532549, 
    -0.093133969274411, -0.0321377731925702, -0.112180372402175, 
    0.0362340659781742, 0.0846452102879683, 0.147633250300693, 
    0.193882081302562, 0.215583612652797, 0.218108100659569, 
    0.184097080705983, 0.157263917364051, 0.224054500294538, 
    0.234981924180617, 0.126698035751276, 0.0843823808665903, 
    0.0959573957727952, 0.112371492296313, 0.117222228544459, 
    0.0894902982934383, 0.0931516811859225, 0.130257347233342, 
    0.129194468291669, 0.0683561700403353, 0.0107319118625428, 
    0.145115022033979, 0.292804298306334, 0.153469810642417, 
    -0.0178218761204385, 0.318556680428706, 0.289168005588379, 
    0.0531375518836861, -0.0390733378250726, -0.162897387734685, 
    0.28503443275432, 0.405784411931218, 0.466554729592975, 0.11625399822937, 
    -0.151525189489218, -0.316957172399794, 0.475421149621974, 
    0.337386369875646, 0.378265812669303, 0.436364405728441, 
    -0.19723242552977, -0.22988856511299, -0.163231566136836, 
    -0.248947447769742, -0.0405776737074214, -0.180271820721425, 
    0.119933962329234, -0.221995690726882, 0.0199900668057654, 
    -0.238332760197396, -0.1999729425518, 0.0376570830614918, 
    -0.144618826170959, 0.0451065101775882, -0.53979303499702, 
    -0.085228580844802, -0.0365220182938037, -0.0424388359117756, 
    0.121582498208808, -0.398280602352066, -0.012155471557613, 
    -0.0615753330492084, -0.0341068817331969, -0.0277854576339269, 
    -0.0269538370568502, -0.0246221740616427, -0.0216930472814366, 
    -0.0168075984740522, -0.0200909503468872, 0.184605522167642, 
    -0.258382397070165, 0.440790447357928, 0.235182748432217, 
    -0.0665531815310117, 0.204790708078368, 0.450048788706258, 
    0.030090533504587, -0.219329113848912, -0.0390944621051766, 
    0.694437819496893, 0.527225504037896, 0.0512212241284152, 
    -0.0542970769008957, -0.354070480960981, 0.732374894009806, 
    0.294768823844702, -0.0861093883084829, 0.0024608248009981, 
    0.567634772503445, 0.416889902264059, 0.234087242572546, 
    0.278235416233377, 0.0204418602839672, -0.0563824233994224, 
    -0.0533151122246005, -0.139873877390453, 0.167053244547431, 
    -0.0227931175843888, -0.0506578835497648, -0.0331581412693049, 
    0.0465490746896862, 0.0284633161626425, 0.00735209921693637, 
    -0.0364688344996106, 0.0752279987335316, 0.0196284743624382, 
    -0.150164460017387, -0.0262960006560039, -0.0802399558309627, 
    0.0435308887397711, 0.0547491146411539, 0.100780828262505, 
    -0.111602803588192, 0.120085877558957, -0.270152997866199, 
    -0.0256737984838114, -0.157268740658452, -0.100839100296914, 
    -0.0884660399489788, -0.101826006609997, -0.0118365039061085, 
    0.0478225058665038, 0.0459363103659529, 0.0509407790839427, 
    0.0469556314653833, 0.0543613000437622, 0.0447177388719247, 
    0.046610425892161, 0.00982929979716882, -0.00603216966181989, 
    0.0748669330804869, 0.0987498012355464, 0.125289958323623, 
    0.184856811386143, 0.180299543294655, 0.10681905124273, 
    0.134248915529684, 0.308122286542312, 0.162287119773948, 
    -0.110675460663231, 0.187236488671224, 0.511052513281868, 
    0.111120084511531, -0.176884023819692, -0.0180616056461702, 
    0.422595168186268, 0.468723985251475, 0.223245821476243, 
    -0.197910473785621, 0.28288851330377, 0.35580992673712, 
    -0.00202477390873154, 0.442877629321522, 0.470396518048037, 
    0.141071241024713, 0.142932524016467, 0.167141090082687, 
    0.208801406453654, 0.124187030619801, 0.639828754341991, 
    -0.116598103259966, -0.116555037314049, -0.118037218057783, 
    -0.115503595986084, -0.112148049757857, -0.123454513277718, 
    -0.0623872841180887, -0.113429856164317, -0.155786237421371, 
    -0.0850275423095292, -0.0252693775414995, 0.0784251530897539, 
    -0.0505509890284577, 0.0354553925226658, -0.0825290965860657, 
    -0.0345410035696479, 0.00492561895000064, -0.0395270823776729, 
    0.0334928235888596, -0.083241643258351, 0.147762860518164, 
    0.162608316207978, 0.00428087645713428, 0.151905746639888, 
    0.219527176678752, 0.215376679365875, 0.219563347802373, 
    0.0902922727122035, 0.104510301428158, 0.401751393522723, 
    0.354883406581442, 0.162509446232214, 0.0927662624911853, 
    0.086439141618559, -0.0362033724968777, 0.0151143273637077, 
    0.376081051739973, 1.1717764067702, 0.138713972498571, 
    -0.238380343023699, -0.391915364741306, 0.192316077266222, 
    -0.308315760669311, -0.0668312736965697, -0.173263209580961, 
    -0.15948574612256, 0.00422911513481046, -0.0784667473587741, 
    0.171405036186416, -0.172708578110767, 0.0787017879342793, 
    0.119758253960945, 0.142184807807833, 0.131669067823029, 
    0.159641750703857, 0.162605943959332, 0.172966850855645, 
    0.142137295774695, 0.155051311899654, 0.108911717313986, 
    0.100404156761336, 0.0931553643292431, 0.0921832841267352, 
    0.105781405240512, 0.114041353280163, 0.0848648645592867, 
    0.0754888972074331, 0.158374626003609, 0.128520019074243, 
    0.0566705750442894, -0.170434737525591, 0.168848659736954, 
    0.418990343614483, 0.0841628203145206, -0.0802722493948602, 
    0.0349301523165566, 0.499295935228031, 0.0249413349543494, 
    0.0859831769985387, -0.188670819576663, 0.540143878755073, 
    0.306654505950654, 0.361331899365202, 0.237188178065572, 
    -0.232993939317798, -0.0869372022152906, -0.380775984491415, 
    1.07719466470693, 0.115736589882302, 0.203352736756651, 
    -0.32223945377326, 0.192112265228247, -0.285496370081918, 
    -0.0681821655348669, -0.202438802889651, -0.109761039899634, 
    -0.150339098810434, -0.161830735214817, -0.0183416089900171, 
    -0.185801661864412, 0.019678407731671, 0.0803226340557418, 
    0.170831912549015, 0.215139058759928, 0.210801740340308, 
    0.181380990605158, 0.163718274282749, 0.195509209337719, 
    0.219081853956177, 0.193793021226657, 0.167557400415056, 
    0.164072987436831, 0.192247027570764, 0.215786882387917, 
    0.217793082242919, 0.222918431282784, 0.229228047126272, 
    0.21770033067557, 0.214462487455306, 0.239588557857785,
  -0.333571703080534, -0.159813735178593, 0.100696129521882, 
    -0.144734814263078, 0.135668816893813, -0.0447653152062485, 
    0.0850232861769639, -0.0750084664649027, 0.0471294701959631, 
    -0.238072288460694, -0.054578800058942, 0.0194535245905817, 
    0.0777283944985711, -0.11545654457974, 0.132613534006766, 
    0.118738583318635, -0.000787624773187986, 0.124020466844683, 
    0.208447348552922, 0.199464192730389, -0.0364242264975229, 
    -0.241510914970451, 0.398887360290913, 0.905076459953963, 
    -0.0786422535518273, -0.132094640431168, -0.346399268718043, 
    0.641893057262507, 0.38902337986359, 0.30914218250436, 
    0.0390580796558561, -0.205199995261988, -0.103752299346971, 
    0.00130619430911955, 0.202693959612931, 0.179543668977802, 
    0.140308542308876, 0.230678062013026, -0.0154524152083436, 
    0.0513438586763893, -0.300411009094966, -0.0462681735665568, 
    -0.122277342795642, -0.30000176673182, 0.237303774716896, 
    -0.210567006200312, -0.0545841634879019, 0.0436417514213411, 
    0.17917183237755, -0.184404114524717, 0.221635915065462, 
    0.314897559102055, 0.0779984732204504, -0.11046011161831, 
    -0.0617512466063292, 0.401033230587191, 0.133826938763003, 
    0.117813399947232, 0.697405970975042, 0.213251102011874, 
    0.0590077080896199, -0.177818744289024, 0.273060213763313, 
    0.63043631202458, 0.283796203597553, 0.0125201683363506, 
    -0.0825373663214073, 1.03788730460962, 0.171369243098199, 
    0.00571400570737515, -0.205933807653447, -0.00670047656971542, 
    -0.239351463274725, -0.0437457675075162, -0.237502315940961, 
    -0.120795882230337, -0.136425599595508, -0.176832547577357, 
    -0.0284424740337002, -0.175135094988642, 0.0303380936635454, 
    -0.001735420716921, 0.223887906112354, 0.161985246780315, 
    0.020386854358555, 0.30146806164593, 0.241798043037093, 
    0.0704473155853059, -0.275222975595637, 0.0964032751885652, 
    0.556939478146121, 0.033980761844169, -0.481599431859957, 
    0.0741567506192753, 0.679394550101718, 0.138751101080068, 
    0.163158158479118, -0.314826317621935, 0.107575536713114, 
    0.545092205427356, -0.393036260992594, -0.283341474382227, 
    -0.144944824498133, -0.314977637218908, -0.144489115200612, 
    0.0293269199581443, -0.231558295519611, -0.053682230541204, 
    -0.0183894594826473, -0.141741373263362, 0.134281438365971, 
    -0.169935260262495, 0.0979648909987153, -0.00195322281365823, 
    0.129310662801088, -0.187583131565136, 0.0631368507139965, 
    -0.152141353537676, -0.0407464834390999, -0.485677917209421, 
    -0.111033855917787, -0.00948239569344836, -0.00693266377191537, 
    -0.0967968383332816, 0.0912250256926297, 0.07388841098826, 
    -0.0226915707811604, -0.0190636713277845, 0.113270912537826, 
    -0.353584940448985, 0.106636883525502, 0.371232441986108, 
    0.582455901505643, 0.32830066853915, -0.0549623719295389, 
    -0.0976105623342631, 1.05207351375333, 0.238369376080288, 
    0.118676897440382, -0.13631335655679, -0.125237670601347, 
    0.26309811426366, 0.797192731381795, 0.326439786476665, 
    -0.0871919114747594, 0.394670886266663, 0.473297498867506, 
    0.154243014830429, 0.118560244415849, 0.609306646603966, 
    0.163368139101596, 0.0215971691796716, -0.017961209871494, 
    0.025468085580738, -0.144399963635926, 0.29111221202112, 
    0.0330915033006884, -0.0865955502558197, 0.0181252711869348, 
    0.209514688076539, 0.0810537788144467, -0.0184897906791118, 
    0.0933219171708237, 0.207397019136988, 0.128350331826131, 
    0.0589607252275209, -0.00116446419109489, 0.188534611889112, 
    0.144064016518473, 0.046376195217946, -0.133821028885943, 
    0.21438211121615, 0.436513466719064, 0.1112496076643, -0.106488627813884, 
    0.013290374195674, 0.396264109171801, 0.204015183684914, 
    0.175988395476059, 0.17871819293139, -0.348150796256688, 
    0.228461212287753, 0.54946671466458, -0.220045081203269, 
    -0.000139515044511332, -0.164652284719797, 0.489642237239946, 
    0.183268549687839, 0.165429833698709, 0.360784277531596, 
    0.00689328530621801, -0.140289651976058, 0.0843059950562735, 
    -0.173152709291183, 0.0404399555939154, 0.0127241823377331, 
    0.0640740114926042, 0.0640179124382083, -0.0666423381695741, 
    -0.0515360920200767, 0.0504356534020964, -0.114360477702398, 
    0.107522406309746, -0.0589670954374478, 0.0990362441085219, 
    -0.0885719129499991, 0.095891340285321, -0.0533608001752604, 
    0.107554692983156, -0.00132079150388116, 0.245652730459008, 
    0.00635998615842349, 0.102658079060177, 0.358682567224806, 
    0.00210461063782748, -0.00284329091538174, -0.0860128136444985, 
    0.258434130061329, 0.148582996139726, -0.0495018587559969, 
    0.550233954129567, 0.323536678536946, 0.092211531770798, 
    -0.20870146739604, 0.383578840851349, 0.0112762858159381, 
    0.344261356259242, 1.15959159383427, 0.371438243787385, 
    0.0664123771475643, 0.230731969288335, 0.422043368012939, 
    0.247962635527425, 0.162611333698727, -0.104841534341935, 
    -0.0550347737617712, 0.43107081424618, 0.170782469722364, 
    0.0449673277580182, -0.0956964794899791, 0.277990589772342, 
    0.276763763181262, 0.0810568920272563, -0.000332027604273602, 
    -0.15587286231607, 0.0343342081460898, 0.406281834561824, 
    0.16402074973526, 0.0318420969026491, -0.152683686763521, 
    0.00200430066068202, 0.284345630244456, 0.164447222867806, 
    0.227870855929244, 0.368394205136335, 0.127820754648102, 
    -0.04004968374191, 0.637624857485745, 0.13369921986791, 
    -0.0397316932603761, -0.206680776284436, -0.0321783739305824, 
    -0.226662381036911, -0.144499790039367, -0.0932832730898407, 
    -0.20349988386474, -0.0880081556050008, -0.120483091831243, 
    -0.148789961578668, -0.0527907574172813, -0.0498123632215212, 
    0.0103977696569094, 0.0551959823967997, -0.0138045303895168, 
    0.0676164537130808, 0.0220150401755573, 0.0415181220008874, 
    0.0660538749930798, 0.0552050430075979, -0.0256925441861423, 
    0.0436627447640423, 0.0904230155115145, 0.0968873805519876, 
    0.121887997416517, 0.133528129586153, 0.0979748093876182, 
    0.0955056987362251, 0.176245183503859, 0.124761839476281, 
    -0.0218018668598801, 0.237184029589164, 0.255663739246448, 
    0.0256029573118731, 0.335453822071315, 0.431661446017406, 
    0.132479868367971, -0.0697758048324084, 0.24445313068874, 
    0.543310249927307, 0.271165377258365, 0.0510591420126096, 
    -0.160378826321265, -0.136276495062301, 0.608235298070063, 
    0.314473371982158, 0.092667384282727, 0.033353138329938, 
    -0.151294485630261, -0.150669310053165, 0.58757713406945, 
    0.0037464376732675, -0.0752412769577215, 0.0157567471731416, 
    0.195075074856873, 0.0104882413170101, 0.00689938274510742, 
    0.0691595827749564, -0.170251099454754, -0.196086555676045, 
    -0.0333493884528171, -0.155652658456879, -0.167599508950105, 
    0.0739295142921194, -0.0685759891332511, 0.117033950074116, 
    -0.109403025199537, 0.019474297514799, -0.181276197144071, 
    -0.0488129906934267, -0.102881652644633, -0.14371073135177, 
    0.153657875966724, 0.0335840006302981, 0.00616131198839248, 
    0.256804303242444, 0.05584949494323, 0.0427834586997304, 
    0.165203112576539, -0.221608379055495, -0.0227590956116004, 
    0.631471007333676, 0.188938919831359, -0.0916992890086203, 
    0.822116859903349, 0.443763869247531, 0.208861453340393, 
    0.311567597708246, 0.412792907810741, -0.295129150798086, 
    0.725980750748263, 0.269015851547673, -0.0582615510558338, 
    -0.0826390811304173, -0.0791434940962989, -0.0584086727889695, 
    -0.0478236341850697, -0.0437470845216464, -0.100295066318166, 
    -0.101812910341968, 0.0508249948061749,
  -0.133905027345144, -0.0954152583183756, -0.305494757231807, 
    -0.143689769018868, 0.0794105984541066, -0.207982954978126, 
    0.0239183354253479, -0.0334326184146888, 0.00939160891536157, 
    -0.227996822881166, -0.0252522650296427, 0.0305735135003774, 
    0.0557656007815948, 0.072009820253419, 0.0756684786394715, 
    0.0566465272311508, 0.0441578901163504, 0.211597631506083, 
    0.143633854312111, -0.220556739484666, 0.159487035511236, 
    0.370152483692315, 0.0932704623881068, -0.0702800888117941, 
    0.220588609885051, 0.478829814494198, 0.41425943734869, 
    0.206756973972475, -0.0232775000994567, 0.762523787291735, 
    0.270284129163122, -0.0331566668711488, 0.0861336988576427, 
    0.448430912106252, 0.254042156585158, 0.17979318662378, 
    0.169002020067812, -0.0929039077134797, 0.462868391300513, 
    -0.19483082226403, -0.33983388056561, -0.138036434423044, 
    -0.299549751648928, -0.263109525616157, 0.151631110674065, 
    -0.278210202412645, 0.0620613796574608, -0.106732226715658, 
    0.0912402232775418, -0.209159793389248, 0.120362387710931, 
    0.111054128627772, 0.103730318391888, 0.143854254512811, 
    0.158854447427767, 0.0920288543459589, 0.111185407138726, 
    0.167755481856667, 0.122691432985835, 0.052364403480312, 
    0.0817370448947895, 0.113829967613008, 0.114793767377464, 
    0.139649035892242, 0.148226039649493, 0.100738423423981, 
    0.155775091269645, 0.225104682159869, 0.102390469868691, 
    0.074255067734047, 0.231701766928651, -0.0250671368430307, 
    0.381004578431301, 0.621268167446455, -0.182639714412262, 
    -0.305661598184415, 0.086612283891501, 0.561263535346109, 
    0.103288005617331, 0.187806190436646, -0.15400522867062, 
    -0.384797047377002, 0.40750283497211, 0.651417583667711, 
    0.0644601634274355, -0.339559868126363, -0.0472989743299834, 
    0.466407602764573, 0.278071424137323, 0.32286564876915, 
    0.435768599856174, 0.248582039925355, 0.0858302519576747, 
    0.000640734362766723, 0.258043562424075, 0.122047184336298, 
    0.0562832247093457, 0.0763312785248131, -0.172632558211255, 
    0.16045905793334, 0.232512865075158, 0.187262944378057, 
    0.148476131019367, -0.136363793138884, 0.177916022846973, 
    0.283805361567134, 0.173267370332348, 0.162495526758209, 
    0.128919159956585, 0.0174152038107033, -0.0145798965649414, 
    0.273697756281252, 0.424578137759697, 0.204757397442956, 
    -0.000497907375526199, -0.0887560523736239, -0.0050658195702248, 
    -0.0745319114815242, 0.476233124481683, 0.074676237499994, 
    -0.1071662736438, -0.01544040827166, -0.0960107425628892, 
    -0.0260896209189739, -0.250952047278436, -0.0469015483434834, 
    -0.0578830905567634, -0.133047860690449, 0.163131405842357, 
    -0.222189278497105, 0.00681318272535347, 0.0648400228468337, 
    0.104896393951316, 0.15754281723737, 0.188532207033433, 
    0.217263465646513, 0.231485616551699, 0.206736747237793, 
    0.166295606030769, 0.152419644279853, 0.214505131667007, 
    0.256397922614926, 0.286109804690251, 0.291331925852967, 
    0.234628232797811, 0.188379080733352, 0.311298270203766, 
    0.373606565841063, 0.187974265934748, 0.00668603174455527, 
    0.106007366354586, 0.424452278558909, 0.409973352182782, 
    0.144567771633719, -0.0548430253993363, -0.0677208054955802, 
    0.570077008454168, 0.238599038225293, 0.100845383171017, 
    0.0403494719525617, 0.233824240512281, 0.763615831586547, 
    -0.0134217233983379, -0.032455991246331, 0.0144373529309663, 
    0.33594850068288, 0.0320061605050237, 0.845734371698377, 
    0.42632842063466, -0.0329475858367242, -0.114206614111673, 
    -0.00755849863802288, -0.126693039371569, -0.0876099957633523, 
    0.00764192101658186, -0.10177841824625, 0.0213918112783599, 
    -0.0796084862694395, 0.0262850485406901, -0.101712812452878, 
    0.0122694157710278, 0.119413568433705, 0.153100384815253, 
    0.15433872635177, 0.252106777433931, 0.213877965049096, 
    0.0527431090379352, 0.271584187901805, 0.46733974473628, 
    0.138817489632767, -0.0177352640057457, 0.0425994762004652, 
    0.656894453238779, 0.0547129371086779, -0.0619426557026677, 
    -0.121566578519218, 0.509059371269673, 0.339997480582636, 
    0.170291518053345, -0.111508657774824, 0.155083997807473, 
    0.340999733628078, 0.294667941112029, 0.160159638651196, 
    0.148793202491478, 0.519550894589827, 0.0656370454260536, 
    -0.120532620533465, 0.31905413789142, 0.138341073187015, 
    -0.287910833317631, -0.0795308796060888, -0.15259345856618, 
    -0.115048832564518, -0.170803137490249, -0.182815205699569, 
    -0.0536369826634344, -0.191278991451339, -0.0289929693386506, 
    -0.17955272250536, 0.0064776620087502, -0.0665748839527643, 
    0.0602153355919528, 0.0138403438739227, 0.0868494629889921, 
    -0.0781299454551271, 0.0729004104927347, -0.0830586693649566, 
    0.0369021804706305, -0.206278314275364, -0.0289284117392939, 
    0.0127335216213463, 0.0788242797576836, 0.123841013577943, 
    0.0897658547602881, -0.00545367727348964, 0.0892783852210433, 
    0.329394516900532, -0.052755723137344, 0.100862548660209, 
    -0.272196543806091, 0.609822057402285, 0.134402726379854, 
    -0.223572711061016, -0.0272488615005899, 0.635899509427025, 
    0.295334159202539, 0.106569553159742, -0.152048894310375, 
    0.0570119558978389, 0.248336643306294, 0.291223460275174, 
    0.400842428253206, 0.4888464411226, 0.266023972308834, 
    -0.099575186957706, 0.45505859032139, 0.250149602391265, 
    0.241993701518205, 0.373901987275372, -0.0410850212660186, 
    -0.0853341873544129, -0.0814361745739853, -0.0097861380438794, 
    -0.190782044131165, -0.0582415584832674, -0.147790389450363, 
    -0.0714864760018062, -0.0124660851077445, -0.0747304820339629, 
    -0.101873408243363, 0.00413235771584956, -0.027616560860506, 
    0.0108641563775926, -0.171518900141444, 0.00596096624585248, 
    -0.115758811439031, -0.105743661545894, -0.0247064633740728, 
    -0.13890574641644, -0.00364335557586233, -0.0589751082717435, 
    0.149179517577934, 0.225215004780711, 0.111080614737732, 
    -0.0514005036462881, 0.153127357058603, 0.230079586637439, 
    -0.0320918273617558, 0.404338240494755, 0.491752150869459, 
    -0.251058783414247, 0.375226369428169, 0.469906057518845, 
    0.664275602681508, 0.92795932460988, 0.0100151329160244, 
    -0.254920763200478, -0.223765931322892, 0.0424110974952058, 
    0.256966784903847, 0.105683687257533, 0.0655640185306626, 
    -0.102782327677049, 0.16413686053612, 0.0625283048908446, 
    -0.0801854855361609, 0.130914693271406, 0.174649583909088, 
    -0.0188921574071959, -0.121503013940072, 0.057178453324612, 
    -0.0484170781015611, 0.0470264150382683, -0.338678926739162, 
    -0.0188876104393291, -0.16023603292496, -0.212700817032301, 
    0.0722106984152222, -0.21642324837155, -0.0081694273720825, 
    0.0351613291201814, 0.0861393747362858, 0.15598343021134, 
    0.150788233149705, 0.0928827854336871, 0.108856322245514, 
    0.224167002603073, 0.1989956427863, 0.165860595523565, 0.175747541853528, 
    -0.0160077018228629, -0.0628699953786471, 0.471983676505637, 
    0.479138363871799, 0.163392620089582, 0.00973236861005053, 
    -0.124327028686151, -0.0440447378434216, 0.372250058289715, 
    0.716938037687477, 0.35474337358697, -0.0303779310940029, 
    0.55426607448188, 0.419814426362194, 0.256115753559504, 
    0.222673249855908, -0.128381471693058, 0.446671251794441, 
    0.747141673047499, -0.141316880989227, -0.142288807177602, 
    -0.0878530442384318, -0.148535942647462, -0.0346367928294453, 
    -0.217807745869705, -0.0385033134258032, -0.0456827252312618, 
    -0.138388671323793, -0.0562143145191576,
  -0.277974225479136, -0.0506393906077158, -0.19806595936645, 
    -0.063417360139644, -0.267477773532944, -0.0925576560952582, 
    -0.17466229992935, -0.17159441711401, -0.00154500016460549, 
    -0.132432624227445, 0.127044255236433, -0.0616764577985686, 
    0.0473692475837789, -0.00984185042295499, 0.0526928139486718, 
    -0.0737972200788525, 0.0391633106662397, -0.0699084052787954, 
    0.0108673610003355, -0.126037639751231, -0.0230622094944506, 
    0.0332390438408887, 0.0411713906582102, 0.139976220655898, 
    0.0998788844642192, -0.0252279272906304, 0.0660792097304516, 
    0.218700859283442, -0.0756706893400171, -0.0751355911060553, 
    -0.371697572218379, 0.299660954846328, 0.649612912981181, 
    -0.100956444129598, -0.263543733315838, -0.223649672312777, 
    0.704868280487377, 0.0415513029571556, 0.0858737836455478, 
    -0.128072938975011, 0.321028932444085, 0.393625302833468, 
    0.259656166623648, 0.0919392427727163, 0.192554285024548, 
    0.0119079176620955, 0.425340290510857, 0.465242650961417, 
    -0.394901948502662, -0.228145293792447, -0.509311026047208, 
    -0.119725003543039, -0.413142681710059, -0.240108448230998, 
    -0.320986085686297, -0.208537840884344, -0.284788464123312, 
    0.0312395115347822, -0.255442651222614, 0.0360061891938099, 
    -0.267862422072882, -0.102417079562914, 0.106620017418005, 
    -0.0426501533866962, 0.156639338455875, -0.0116683048613495, 
    0.0956226368627416, 0.044180084109744, 0.0263291696452941, 
    -0.160761306528307, -0.0264563457039821, -0.021716386616414, 
    -0.00759488367272959, -0.00147258832218843, -0.00076298241097042, 
    -0.00161258977369769, -0.0157724347826347, -0.0616352647235575, 
    -0.0152151179091356, 0.0135112162088508, -0.278687399974322, 
    0.593609583507735, 0.276675383400871, -0.17367409543284, 
    0.296018044922913, 0.586366180291305, -0.337974282559103, 
    -0.147870199539131, -0.39334985591168, 0.481111871994542, 
    0.364130882407629, 0.155325743365536, 0.0668137143961637, 
    0.171714428873095, 0.138405252686863, 0.0634892811705999, 
    0.1139358326196, 0.185360951977316, 0.118781240605908, 
    0.0363482904170944, -0.05614060761898, -0.0555665989369593, 
    0.0194739675502306, -0.0593001923710906, 0.0099102496199312, 
    -0.0800700394492103, -0.020157825096447, -0.0452778342058604, 
    -0.0243476494703077, -0.0487574844410661, 0.05428983929004, 
    0.0630852973056243, 0.0963748972093762, 0.253903360906222, 
    0.183641198013537, 0.017951762300114, -0.0502252994442199, 
    -0.0140596413197165, 0.409691407573513, 0.226279012815179, 
    0.093481668671158, 0.809813231769555, 0.263074629878458, 
    -0.100649539765689, -0.239770920685118, -0.0466920683439732, 
    0.887907797169884, -0.106490582390668, 0.053816383343253, 
    0.467096403727805, -0.0864351985739166, 0.0793432804890477, 
    -0.104918918203637, 0.117040145004259, -0.0767918554820626, 
    0.0919161981808998, -0.0542905301127327, 0.0145528654379926, 
    -0.166442808837695, -0.130334800654064, 0.0386640456292722, 
    0.180041762010824, 0.131250503067519, 0.0818054604639517, 
    0.276295592958455, 0.319979094428419, 0.213482302370788, 
    0.203851812334345, 0.285137945150127, 0.229971344753232, 
    0.0807691256372708, 0.0622305633227342, 0.0872351465836137, 
    0.073804421371276, 0.0804766258460804, 0.0464843931392246, 
    0.0585139419807677, 0.081004291266219, 0.0864541202609981, 
    0.0272927633077199, 0.0628442403569168, 0.0810476979477571, 
    0.0891669925718545, 0.107150140467529, 0.100979035426672, 
    0.0777795091119667, 0.0983602133763435, 0.123901288375866, 
    0.173213924817734, 0.132224190253727, -0.115508031898397, 
    -0.012505812720864, 0.526237700613652, 0.29779557623157, 
    -0.00397450306452902, 0.634859276150522, 0.375126155159723, 
    -0.122370326792811, 0.0698108468475194, 0.0986536562426784, 
    0.620752167351353, -0.270549401585089, -0.248681862135302, 
    -0.383173701390081, 0.738218600308415, 0.375855959012708, 
    -0.262551289460377, 0.758829490370864, 0.379967318175124, 
    -0.323894993959034, -0.205310177219688, -0.102392623015185, 
    -0.111359089613214, -0.13122827934402, -0.0435911508809226, 
    -0.136112301292663, -0.117401795131718, -0.163330069813038, 
    -0.116194777222817, -0.111850006888338, 0.118202312895315, 
    0.0631628705749005, 0.0592136046437125, 0.143368041383837, 
    0.164425836826779, 0.107977362165956, 0.0771254623462103, 
    0.168581689400873, 0.181256768786493, 0.127115545520782, 
    0.0753736356392906, 0.087520170975452, 0.0673226912465414, 
    0.0736969334765233, 0.0658002376373528, 0.0649246021465049, 
    0.0661357399932253, 0.057797238149267, 0.068619020229663, 
    0.0608952260268511, 0.0742728355754492, 0.0798376103189123, 
    0.0879515599793702, 0.0734902696579909, 0.0769088109650024, 
    0.0710068457737903, 0.0764278480975371, 0.0959548944291933, 
    0.0868675617157552, 0.0213422278083527, 0.151873572240748, 
    0.173476447156675, 0.0602864592068443, 0.108876603141866, 
    0.342629540681078, 0.244439756401024, 0.102150776646388, 
    -0.044346699346923, 0.408681126551186, 0.235123335733187, 
    0.112840532012003, -0.244563277962425, 0.329549324475976, 
    0.513122360173158, 0.146429151828689, 0.0216202146185206, 
    -0.153732434710542, 0.0530994567453449, 0.306214234759469, 
    0.469548081789546, 0.420502822596028, 0.150724414229763, 
    -0.128404000533534, 0.152081427592275, 0.33274065697889, 
    0.0704403264566028, -0.163591382115813, 0.245608695582762, 
    0.148309022014394, 0.000297875064118804, -0.09784795234312, 
    0.00872093953744783, -0.430809449925618, -0.110309587254902, 
    -0.0349968392471707, -0.280392093150474, 0.0460189256819279, 
    -0.0448645955102812, 0.0732701307301151, -0.262481258388198, 
    0.0136565816062625, 0.0577803053701534, 0.0791649043968875, 
    0.0929336859618696, 0.0962584535281676, 0.0705976875026647, 
    0.0849549997683986, 0.113481011057547, 0.082014540385306, 
    0.0212628628095116, 0.0639173748907757, 0.146426366901319, 
    0.179333829275378, 0.145095419255948, 0.108092139864672, 
    0.167399292273897, 0.29960117238798, 0.192381921872294, 
    0.0179465721879434, 0.269566690499297, 0.352087449334984, 
    0.300886343020268, 0.395008109210685, -0.355589569759627, 
    0.474374982025804, 0.526890979659771, 0.182572101234803, 
    0.573439749136929, 0.580307110420362, 0.161946942143242, 
    -0.0561684463491735, 0.276639906396397, 0.248230404869848, 
    0.0979969309091778, 0.0178225086122838, 0.037375076208268, 
    -0.218045587990696, 0.15164376194109, 0.269591413335861, 
    0.0332438653973527, -0.128703581921282, 0.0884250173461308, 
    -0.149524632308096, 0.0209250653292288, -0.33300192951618, 
    -0.0862118742505739, -0.0992586326928559, -0.23850510251742, 
    0.268231518000169, -0.191539670089645, 0.126025187680959, 
    0.0373533755459243, 0.0450315039879528, 0.0947195853330328, 
    0.0476279830121438, 0.059193615921819, 0.0373628675959799, 
    0.087062867124959, 0.125806014994683, 0.0516824793576829, 
    0.104126883627122, 0.13327636275273, 0.125149466590796, 
    0.187110072602668, 0.221182142289322, 0.131737847355476, 
    0.0864767016372875, 0.269927559991656, 0.31975707636916, 
    0.137100686594896, -0.158602117403081, 0.170423963534188, 
    0.464021806174686, 0.147557160802782, 0.0826589625256853, 
    -0.280971112463102, 0.176484232360086, 0.481060713734193, 
    0.153984636114303, 0.0512386540825143, -0.237015252910556, 
    0.101793605500637, 0.41945377259021, 0.103997980100782, 
    0.0139261996242608, 0.152069835984378, -0.218377335064873, 
    0.397754909026226, 0.41202463636085, -0.289016342927369,
  0.143244706268878, 0.297897972662245, 0.231572329576795, 0.071037635805378, 
    0.120152770765466, 0.521750589963146, 0.21133394020092, 
    -0.202448145200925, 0.415347358092686, 0.332403437949176, 
    -0.136503574124648, -0.192551989407917, 0.532693777796686, 
    0.667567686327122, 0.369462717012498, -0.242278638216588, 
    0.406291444247405, 0.443280473085296, 0.00793306084095605, 
    0.336948226195445, 0.591919547930377, 0.301141155053443, 
    0.138633929741814, 0.0972072088843808, 0.0911994905707724, 
    0.0888998595967577, 0.0940908057287925, 0.103309861576401, 
    0.0909063813322947, 0.0728519279352974, 0.119575279301151, 
    0.125374043008297, 0.0966799216604608, 0.123937122545176, 
    0.173930246232972, 0.125027508373802, 0.105312583736998, 
    0.222913308012168, 0.150283468640604, -0.12916165530732, 
    0.302004971326027, 0.420432094916144, 0.0422932545192991, 
    -0.135141076816822, -0.125543405449455, 0.410137442375709, 
    0.308700175234456, 0.343531890097091, 0.241100025616239, 
    -0.260816109136181, 0.14422703708857, 0.527475507065411, 
    -0.0477637263492789, -0.260103001157351, 0.0996415391817911, 
    0.220143717066753, -0.0851632815430713, 0.893433161531648, 
    0.384771520743597, -0.0314397456988618, -0.2150370550304, 
    0.102643161823582, -0.0782545022693922, 0.0892334199321758, 
    -0.124920042437269, 0.0516851318491444, -0.409328668774725, 
    -0.0763901831480672, -0.148888694067046, -0.224471653497245, 
    -0.0128208353691797, 0.0631783935630709, 0.167978305955274, 
    0.202685514062978, 0.206645748582853, 0.167570675436076, 
    0.154542781651705, 0.227540388485297, 0.250578031632597, 
    0.222797169215342, 0.233476457569772, 0.202123917179249, 
    0.215227973809515, 0.293241360677251, 0.274931878606451, 
    0.222314152729131, 0.27271106911233, 0.22421467641474, 
    0.0881500582459139, 0.496485611981161, 0.392189289160095, 
    -0.0445800164605486, 0.59079278696631, 0.533658851687498, 
    -0.243754224173134, 0.037854270512543, 0.574719851885406, 
    0.320701487170042, 0.484154622561976, 0.440154615730445, 
    -0.245138891938675, -0.179170244515616, -0.151463628723208, 
    -0.239714382875985, -0.0826085597209261, -0.252073376101925, 
    -0.122864037759431, -0.135365972455195, -0.0965670002312668, 
    0.0500540575573339, -0.021691251914562, 0.154633758565392, 
    -0.166296023500064, 0.0350197789229587, 0.125906756808697, 
    -0.23254680710674, 0.0040097891965393, -0.0529872705386139, 
    -0.168632566721491, 0.17586246680813, -0.218661543546862, 
    -0.0702173643835702, -0.042982075665279, -0.0825926913210368, 
    -0.0957966473839618, 0.0086775294846393, -0.0883954902164818, 
    -0.0112360427576409, 0.00588872695372045, 0.106827078574592, 
    -0.423774605509387, 0.882052224277125, 0.200843498501151, 
    0.0423204606522049, -0.20201297669091, 0.804979842222813, 
    0.153291227070051, -0.183384052920421, -0.0100782565300316, 
    0.603067717817017, 0.389744670299178, 0.240459316194461, 
    0.246234467608208, 0.137130014079552, -0.342554151181316, 
    -0.0837271988386878, 0.656070964198926, 0.284038523214065, 
    0.042582846391287, 0.577007428859849, 0.451261161496213, 
    0.155318752850047, 0.0563703882988497, -0.0764748867231952, 
    0.0543606098895274, 0.144702523925893, 0.236522038604886, 
    0.55829765803123, 0.12223722536188, -0.118483205511765, 
    -0.225559574455749, 0.228517671257414, 0.550836849198827, 
    0.150901958592389, -0.132508859130702, 0.000207223828436617, 
    0.186442624201741, 0.76804299625725, -0.109358159792591, 
    -0.234053780216019, -0.362880029585049, 0.0844335629310812, 
    -0.287676995189103, -0.0754280417984889, -0.222914665045734, 
    -0.161984764705931, -0.037085763935378, -0.184136266793613, 
    0.0427292971845514, -0.219479201393766, 0.0203829242186539, 
    0.00322257282903651, 0.0346368712804276, 0.0187461952204034, 
    0.0544098051985718, -0.0679099707811737, 0.0109872310608826, 
    0.0336636419339029, 0.0559237092101939, -0.113293232757089, 
    0.0300729649899616, 0.0315219152546144, 0.0295609643416421, 
    0.0642595921354652, 0.0540928325073485, 0.0316490403798539, 
    0.0299644713485306, 0.0628817701889211, 0.0493888920018039, 
    -0.0040891444416942, 0.0799600123137492, 0.12190883403544, 
    0.120001529256755, 0.149722802310611, 0.208085288502794, 
    0.205082201289783, 0.170850916437234, 0.135306434567442, 
    0.146154387035461, 0.341767940608857, 0.266811661772039, 
    0.00743413577316887, 0.0432403075030246, 0.569531104143808, 
    0.2170481902648, 0.116097619019015, -0.164902118104439, 
    0.576465373784066, 0.229799767548707, -0.0915076326583518, 
    0.338336679298093, 0.433933698551585, 0.183064069391615, 
    -0.231070117791976, 0.547848547520558, 0.353513607761767, 
    0.0676116263636263, -0.105636466200559, -0.0741555913632911, 
    0.542449805484822, 0.184051007903982, 0.0349633010795547, 
    0.29525089413641, 0.175162571055748, -0.166785656997089, 
    0.155850774523439, 0.205588745494247, -0.0992428438054446, 
    -0.0236805760158659, -0.0338712493321901, 0.0280751362089581, 
    -0.22965877725637, 0.0732270569596861, -0.104167066020742, 
    0.0479663522885542, -0.222014070819742, 0.0462883249840708, 
    -0.148680427445036, -0.000574416570683189, -0.237073794299835, 
    -0.0999425475390965, 0.11253978811874, 0.136135645220421, 
    0.0698678562944459, 0.0706494287191358, 0.151066064479386, 
    0.280285367267315, 0.300344234728981, 0.155738335005886, 
    0.00186416372236615, 0.398018221131234, 0.362869932025074, 
    0.0554719037333136, 0.510432232335025, 0.602357374064709, 
    0.103908730200648, 0.174994534257776, 0.92810731115751, 
    0.206390717806853, -0.0772079051578069, 0.195603115490023, 
    0.660042004605826, -0.0914810975790093, -0.0262945283749606, 
    -0.114723334628288, 0.514040239797497, 0.241998819901582, 
    0.0823608936139027, 0.22357032131213, 0.561749291231554, 
    0.0460294915583414, -0.00166548125999139, 0.00925260111066699, 
    -0.114956770529889, 0.180444461972306, 0.0566074668329923, 
    -0.0275358726352594, 0.031514441260797, 0.202186045318364, 
    -0.00619759161749565, 0.00214983762149812, 0.0558094877383074, 
    -0.00380800627177338, 0.0334789797174476, -0.0225206930698294, 
    0.00563011113711559, -0.0171816353393603, 0.0493675424356709, 
    0.166410896717339, -0.227698600274195, -0.0320575671754205, 
    0.410325836533787, 0.439946515191309, 0.174163727779044, 
    0.102163510209705, -0.244101858478031, 0.434759789219569, 
    0.384614416383496, 0.235613898902602, -0.0877398524874111, 
    0.5237678560355, 0.370522252494583, 0.29101344462788, 0.767542908697308, 
    0.446596983084627, -0.29377656190722, 0.568643540496412, 
    0.505537810204679, 0.537702013827979, 0.630640514166403, 
    0.0323753509913857, -0.122042055031263, 0.10983448666199, 
    -0.104760004113662, 0.267790134782669, 0.0841503082635925, 
    0.00797227289092396, -0.0391520421697297, -0.111356059062547, 
    -0.000868001352372125, 0.357248486488861, 0.236508822996413, 
    0.162802426376586, 0.201299620889499, 0.0423600619520472, 
    -0.149649519304164, 0.304634797078967, 0.436807864924182, 
    -0.0948783246557831, -0.140534734676287, -0.231138805548525, 
    -0.0397936804875988, -0.0644021083277799, -0.140608636024338, 
    0.0584012690604577, -0.117786017178503, 0.047715024664324, 
    -0.0346409998455266, 0.0942031793355804, -0.122186848629364, 
    0.0526289625958014, 0.102915564441148, 0.101345797244769, 
    0.138654579297825, 0.15885710214713, 0.128096672274723, 
    0.121760174692512, 0.158689264518294, 0.134442584910722, 
    0.0545414549718609,
  0.415442902622747, 0.0401768285358671, -0.223625720130993, 
    -0.0594702134960646, 0.417770047001953, 0.358220480783468, 
    0.124796022954105, 0.036508954517087, -0.228414248134239, 
    0.322668123248958, 0.393792592088779, 0.153161084017361, 
    -0.00937252008322492, 0.391202923337174, 0.326082681127367, 
    0.0719786040863669, -0.0695156047838357, 0.0652420329759033, 
    0.457538036152171, 0.517547656780323, 0.133420518056047, 
    -0.143390115594817, 0.142920063218704, 0.304885202678227, 
    0.0476814632818253, 0.0406481787884474, 0.377690543655048, 
    0.217474376705042, 0.220790979106025, 0.39735698768576, 
    0.107308609450608, 0.00317258383863162, -0.0107910402093221, 
    -0.0869896835844015, 0.00814316849998092, 0.0157841191406611, 
    -0.0719361747499306, -0.0650496705557985, -0.00245777930125696, 
    -0.00568545740158855, -0.04456778147537, -0.0575076743624997, 
    0.0455874236090896, -0.0178296764792752, 0.0405983414874571, 
    -0.195227332772956, -0.00802888458069402, -0.062164626111209, 
    -0.00812179002024474, -0.247676481848612, -0.0658801895119985, 
    0.0977723481443092, 0.036856497298628, -0.0328371253439552, 
    0.150494231254245, 0.170867073411309, 0.101246679811895, 
    0.054835335559539, -0.0290756960370171, 0.0757020811440626, 
    0.672777498850532, -0.0413407705716829, 0.077326724917435, 
    -0.20486380333655, 0.326535765964702, 0.315569643300657, 
    0.683758384460506, 0.344880373408063, -0.147803329135312, 
    0.0185055629192875, 0.471086148411214, 0.226665701717337, 
    0.289461109521475, 0.225027588169752, -0.0571441722719991, 
    0.321070226953419, -0.138648651787035, 0.700716200276729, 
    0.178322913320558, -0.160144632608242, -0.208699925926317, 
    -0.0733331076102987, -0.122151904746073, 0.00340157331200656, 
    -0.201373444242566, -0.139677455829406, -0.0766048892968088, 
    -0.233290521942529, -0.0881070264819909, -0.0651692159182517, 
    -0.188557337404828, -0.0636632283805599, -0.16058629897879, 
    -0.0377329312437072, -0.0792788737718997, 0.101480473408472, 
    -0.0121175300361086, 0.0657234777042334, -0.449848882198258, 
    -0.0847747612665674, -0.0278784348695335, 0.00799668840849643, 
    0.0836961098486488, 0.162947343683697, 0.129381319087818, 
    0.0907818115804126, 0.120889303698925, 0.138519559944329, 
    0.142096609886638, 0.161769690854795, 0.215093819689727, 
    0.206855382390308, 0.19827108432695, 0.221599765916418, 
    0.223362236831248, 0.14524344393053, 0.124955905136843, 
    0.386161464761383, 0.235427924399365, -0.0843857376650776, 
    0.186793812542821, 0.478623120351973, 0.328585543862977, 
    0.0964293979841725, 0.00280793762095045, -0.295886582150304, 
    0.540170815709769, 0.282728543293293, 0.140243420302651, 
    0.0585773847111965, 0.107955824002511, 0.198222471401589, 
    0.0773596430387343, 0.0151100256221687, 0.27194276316552, 
    -0.0350108490013628, -0.166099573726746, 0.0459439319967485, 
    0.188483233377724, -0.102247550085187, -0.0242194380979408, 
    -0.222202088709406, 0.0437908886790208, -0.115642229114049, 
    0.0152727209775244, -0.240760216474972, -0.0129168976304024, 
    -0.195283512515279, -0.133100865842973, -0.0707662881103724, 
    -0.202997603913312, 0.139345124236903, 0.104668838204431, 
    -0.0195610824247193, -0.000601056813392786, -0.0486780796892667, 
    0.3903142812286, 0.110048953602706, -0.122292525502988, 
    -0.00275432403084067, -0.491514835890578, 0.271967392194688, 
    0.608754926333381, 0.602599149795642, 0.153673330452863, 
    -0.302888306155997, -0.251804679954967, 0.721875475304512, 
    0.316258121673105, 0.00126360256075528, 0.25476937106909, 
    0.38053557452734, 0.0560496115486642, -0.0510700164949012, 
    0.0350175241691438, 0.340255878775387, 0.570315735574165, 
    0.307179356140987, 0.127963060147536, 0.262544101847822, 
    0.0879544486416287, 0.147509232633993, 0.303456656411611, 
    0.088997963093222, 0.0212597171864196, 0.0490304988719423, 
    -0.0336397356166687, -0.0228012915763861, 0.330328874732245, 
    -0.0304595036377281, -0.0337897705470583, -0.0141361584371588, 
    0.043638679214233, -0.0529084162598392, 0.0283775403159873, 
    -0.0371038474667652, 0.0475720717959585, -0.0232853486824783, 
    -0.00877876533894142, -0.0315421236458018, 0.00957723971935753, 
    -0.112401147670625, 0.039583041594112, -0.0654584501467599, 
    0.0159760814590468, -0.130525457132168, -0.00992417486769914, 
    -0.0851803036230472, -0.075743440076905, 0.0181858804506883, 
    -0.0752422442043322, 0.0364793639700904, 0.192261431303041, 
    0.156999574530035, 0.103877983455153, -0.200171265223382, 
    0.209712629929069, 0.381045624709916, -0.0172363736140397, 
    0.144449511030542, -0.0129240860044926, 0.575722445239161, 
    0.174785486922513, -0.158508248874687, -0.0503264425241022, 
    1.31724255299497, -0.0863825396589999, -0.369621668164718, 
    0.192570081694014, 0.617530461786957, -0.0919383368200989, 
    -0.093240663577568, -0.0898840374788181, 0.36837972610609, 
    0.182342400009233, 0.040723491779928, -0.121752807027285, 
    0.118997715596728, 0.303711983342866, 0.224687740308065, 
    0.139725581927237, 0.127596919863998, 0.111486648512296, 
    0.0979297082537543, -0.017873923768561, -0.067698173276681, 
    -0.112506553051407, 0.101546518768927, 0.0851100325532608, 
    0.0225372191748434, -0.023704156890118, 0.0589992423063431, 
    0.201832910070971, 0.193474605944884, 0.108976047279843, 
    0.0265333001139856, 0.056102719313127, 0.195909781100425, 
    0.16715172385581, 0.0793615890872388, 0.0103217658121973, 
    -0.00680931538870451, 0.0220880725758099, 0.0315216029399084, 
    0.0483114148542053, 0.0170125811919251, 0.0623144788100699, 
    0.0487006582313843, 0.114226621997328, -0.086119459761845, 
    0.150442467683837, 0.279212593008019, 0.222166333104512, 
    0.136457318881519, -0.131504508010399, 0.290290802879072, 
    0.384387336532269, 0.29119892110136, 0.118345400605672, 
    -0.243449927170129, -0.104651377745272, 0.890277814616979, 
    -0.0122756163460307, -0.276452970751565, -0.221750246144495, 
    0.689762199575551, 0.324188928040408, -0.0634297702138773, 
    0.697839282296406, 0.318066547260591, -0.259079226372505, 
    -0.0700904565023329, -0.148510016247282, -0.045877157962948, 
    -0.0955697347908557, 0.0704724570358089, -0.248523467829517, 
    0.0952985398261021, -0.159801135898215, 0.216989397794601, 
    -0.0983055571442309, 0.216450624210731, -0.162558535447068, 
    0.16614058728348, -0.105739701764892, 0.158927719362516, 
    -0.249233053156047, 0.0508032748101967, -0.241333161581904, 
    -0.10290342484929, -0.0499156669717286, 0.043136144565106, 
    0.0301808198470702, 0.041456530081028, 0.00714136539133276, 
    0.0214970389716832, 0.0114988371066086, 0.0401413351070918, 
    0.108157233906374, -0.140436349565927, 0.267581820636929, 
    0.250173074273363, 0.0964030838488506, 0.286938536549497, 
    0.247242143563662, 0.00896936575382146, 0.370756956133741, 
    0.686382786857283, 0.205017248811735, -0.353819348222711, 
    0.239843067512154, 0.445752183505783, 0.98073996830425, 
    0.733448636419433, -0.369819640122408, 0.592075460128229, 
    0.451688916389495, 0.598941780618513, 1.04557078199459, 
    0.00910847695812193, -0.203324796942279, 0.104499021588387, 
    -0.186472937693932, 0.22758019071468, 0.174870359724135, 
    0.0249093584434547, -0.0347535987646382, -0.121592512549741, 
    0.282278424269688, 0.0436321338091324, -0.0103930980745752, 
    -0.0199596723971857, 0.247899511427929, 0.0630310291057546, 
    -0.0490136697367195, 0.10113718412764, 0.189444760741394, 
    -0.0798733635214086, -0.103169513255956, -0.106959895114548,
  -0.388213090854816, -0.21130769259045, -0.175125871100806, 
    -0.12608490536477, -0.154876599978109, -0.168601161326634, 
    -0.111757679062526, -0.289313053042425, -0.0711121295774639, 
    -0.183676467308225, -0.0215023623014448, -0.0312633211464163, 
    -0.0620423351082941, 0.0221164980755373, -0.0850961924771772, 
    -0.0115430549453453, -0.00334979380741506, -0.0303225919943036, 
    0.0787562998979158, -0.0709600930083395, 0.0216871369849706, 
    0.0679254234495805, 0.106658721543711, 0.133482880506943, 
    0.13517388963998, 0.131491296362567, 0.1434595413919, 0.15573529831286, 
    0.133603453460789, 0.113312405360189, 0.149779470154362, 
    0.15860492795172, 0.174351487576355, 0.222316197708579, 
    0.250968944742341, 0.193873746922104, 0.108658119282691, 
    0.193390938876683, 0.337830116134105, 0.171172908753707, 
    0.0477256916650381, -0.0919449619083979, 0.361339146832583, 
    0.466107613699279, 0.18705692692796, -0.186271073167679, 
    0.229777102074749, 0.465246650808242, 0.0867695377467801, 
    -0.292507522055596, 0.0458860533519927, 0.578538357396705, 
    0.304650662653765, 0.18917790979703, 0.200345482510754, 
    -0.045211082336977, -0.175845066780743, 0.21628897956372, 
    0.860741592956338, -0.242882316583711, -0.362424763366004, 
    -0.145995776090152, -0.190221387654897, -0.18011658309053, 
    -0.179271881365254, -0.169426921290617, -0.104001794029873, 
    -0.170246529920427, 0.0663352684938685, -0.229186706497392, 
    0.116000619102175, 0.0123314864930529, 0.0493312389213756, 
    0.0577020895167483, 0.0746985712453917, 0.0114345325957801, 
    0.0598859449865994, 0.0486181544261836, 0.0748669207961642, 
    -0.021083715891255, 0.0428214401102282, 0.0489538069707399, 
    0.0434011807627016, 0.0130222829533374, 0.0414258917212932, 
    0.0214558348724878, 0.017777898554357, 0.056987792559097, 
    0.061590915033266, -0.0316305239267686, 0.0495736547328587, 
    0.190332490407593, 0.133364538059737, 0.041052040982402, 
    0.150895714478704, 0.285802832686699, 0.161758541350523, 
    0.023841317536883, 0.41579839697476, 0.238035248561413, 
    -0.169237973020861, 0.0540698126929128, 0.664828252406313, 
    0.130953298607664, -0.124320674423769, 0.2940262985354, 
    -0.107112426907968, 0.634186055102642, 0.769915756004622, 
    -0.0375581429071039, -0.152060525297199, -0.114206829802274, 
    -0.00671326097401566, -0.00814942354077153, 0.0310656919389411, 
    -0.161891030207671, -0.179616403644775, -0.00119915509773641, 
    -0.20287522799782, -0.134368073124633, 0.118104775006858, 
    -0.266034997540632, 0.110551524929116, 0.0686719608265245, 
    0.152206131576305, -0.336843899179005, 0.226578807138312, 
    -0.252313678255134, 0.0607403043662427, -0.251629979970577, 
    0.044731887357379, 0.0349222545395527, 0.109245007671022, 
    0.151559692464811, 0.13949109972641, 0.126318084521293, 
    0.101701624677568, 0.137753897396257, 0.165219919248834, 
    0.156232429456441, 0.162504613251828, 0.129388147348247, 
    0.122376255294945, 0.12579076298048, 0.17044530468181, 0.136459750076042, 
    -0.00576900037394129, 0.233757086136065, 0.216246416269353, 
    0.136516737929442, 0.292156102060195, -0.2371292961135, 
    0.272635015748951, 0.625259283987793, 0.176842042733841, 
    0.101297861184073, -0.00125625019674583, 0.248129510411393, 
    -0.148982481501925, 0.241965457469029, 0.843602653224281, 
    0.286415743207994, -0.084103987405214, 0.669117298801426, 
    0.364858528197689, -0.0178921975081896, 0.566191604616319, 
    0.50706463603358, 0.126487824670811, 0.44430639040952, 0.389454606718091, 
    0.0605967624914571, 0.0124136802763566, 0.00566189428355105, 
    0.00833280014195267, 0.0427285361036848, -0.0510843669904685, 
    0.100684516651111, 0.041536022477697, -0.0847590024332165, 
    0.0593408142374736, -0.282706515999533, 0.246352208370542, 
    0.518517537658789, 0.0914441908634651, 0.00250691463996855, 
    -0.255607468755319, 0.323978740168541, 0.425863707656918, 
    0.141154686623738, -0.103862110744994, 0.0857595326431304, 
    0.404600128471175, 0.177347108824995, 0.0368504847051585, 
    0.174983739979175, 0.139926945773986, 0.0540325888265681, 
    0.516891917974555, 0.24121383120293, -0.0254634646236629, 
    -0.00973711117401724, -0.0248979367124352, -0.00732457881055487, 
    -0.0218802011114296, -0.010127315650412, -0.023952985114822, 
    0.00259622482432315, 0.0576314686168145, -0.112267850932063, 
    0.0862817908687625, 0.181273170678829, 0.0253812850731848, 
    0.257087366045144, 0.303032545776147, 0.119132368158847, 
    0.012932482005556, 0.0934955473978035, 0.529784354088771, 
    0.186899480210693, 0.0609716630895116, 0.143233066246075, 
    -0.0656158990907613, 0.108918970251298, 1.03807914137184, 
    0.0759623205047564, -0.0417694578839994, -0.118766335365628, 
    0.749034262806024, 0.137381117170558, -0.046717945066714, 
    0.0485008453384297, -0.0566716274441018, 0.0265515636715431, 
    -0.0750623509845417, -0.00650805410952952, -0.143379415190087, 
    -0.0505608195889728, -0.0428820810818728, -0.0853955021169777, 
    -0.0219004007558048, 0.0888511001693923, 0.1667781490642, 
    0.177628281720349, 0.172361708100482, 0.145444214235387, 0.1925607459515, 
    0.299322938035841, 0.235100945945021, 0.111521700793934, 
    0.127090106024967, 0.344056889203986, 0.328171680712564, 0.1587167078699, 
    0.0732289969340913, 0.140996457782896, 0.387424467444103, 
    0.554730819239559, 0.197691078180877, -0.117650085753772, 
    0.000467691340274551, 0.614544853388439, 0.249486520853887, 
    0.177944593499299, -0.222883112679019, 0.259776491709989, 
    0.467791515806044, 0.234324245770071, 0.0387123019736399, 
    0.128151348570597, 0.107271209210606, 0.244653556120524, 
    0.184124684779824, -0.025370303175089, -0.147737243558338, 
    -0.00467688451825859, 0.0879390156814199, 0.0818798058143656, 
    0.0136947572823393, -0.0563520225153443, 0.0152960529436535, 
    -0.254113554511333, 0.0540846587814152, 0.00263825174952156, 
    0.118969320442029, -0.212504111773041, 0.059538792065918, 
    0.0382780708583476, 0.174411367615212, -0.269856999645805, 
    0.125083893799604, 0.0843876808074266, -0.0175328527690052, 
    0.0466114659574811, 0.310091401090063, 0.27368662737102, 
    0.156641074541174, 0.145834123088301, 0.155422106842995, 
    0.0572514602945312, 0.173366461714676, 0.428986982400512, 
    0.455781165151661, 0.315142377766846, 0.451920168949445, 
    0.745117322257235, 0.443705229760936, 0.0908756473141553, 
    -0.0167193010978924, 0.786325061092049, 0.450721295262787, 
    0.0866660305074263, -0.368384924705817, 0.003419299035419, 
    0.519624270510781, 0.28822134472566, 0.24601661558551, 
    -0.280754653044836, 0.46436560222057, 0.323262936254807, 
    -0.0214973815375636, -0.0526315379439212, 0.129884147473056, 
    0.147828964664112, -0.140380247286895, 0.274188788099649, 
    0.0564496393242494, -0.092474935031672, 0.00226776798384891, 
    0.254161234851662, 0.0597385443255428, 0.0179267563793074, 
    0.0103955735887337, 0.00838575838741548, 0.0188699461224442, 
    0.0124331804124323, 0.0129322061705066, 0.0212367120557921, 
    0.00124936638995873, 0.0148341513532371, 0.233763960213726, 
    0.115126582048054, -0.0725312593954055, 0.264358751288182, 
    0.26070186024558, 0.0590028046100698, 0.295321312878862, 
    0.474011430086461, 0.350385389436673, 0.227516645069284, 
    0.133332324551166, 0.0260074500645502, -0.217057223025805, 
    0.0852852646690807, 0.31595306243376, 0.178968129754701, 
    0.317417790890089, 0.755691301467329, 0.867418525958931, 0.133838338260454,
  0.821280449743619, 0.25324524869399, -0.255133324601151, 0.461961036175794, 
    0.42164353573737, -0.0924259645335632, 0.321473500231951, 
    0.0721267033490893, 0.71658628916128, 0.0444966994014965, 
    -0.0861031287976529, 0.0609713891466364, -0.183167182256151, 
    -0.0385037970805346, -0.0372686768571651, -0.106383605022036, 
    0.0502478689064315, -0.0240729379345089, 0.083677134346779, 
    -0.12017787072786, 0.0366556419180556, 0.0926874505655161, 
    0.126723033476618, 0.1876291786729, 0.248706207828094, 0.23898946089552, 
    0.209716022138832, 0.223300419147067, 0.227420485965853, 
    0.23266442931681, 0.311282905911591, 0.280702186437751, 
    0.173345534768362, 0.236658551796134, 0.458858400726113, 
    0.316075728546416, 0.0973316426634929, 0.0156481499001231, 
    0.453479257577136, 0.490103930351566, 0.141283775319718, 
    -0.162854493820501, 0.0602469053004193, 0.56131453472418, 
    0.234852920915036, 0.136752928592635, -0.104410566326922, 0.537679010432, 
    0.235919072312163, 0.0512799218056753, 0.283106084283718, 
    0.443257327481637, 0.263547988146586, -0.243411827404205, 
    0.641980520527268, 0.144830040428678, -0.0713386927244691, 
    -0.0169425197006162, 0.0919137810663013, -0.10032925806229, 
    0.337806194572219, -0.138571607080413, -0.209126962765723, 
    -0.264528249211883, 0.0218842907360891, -0.133905402698292, 
    -0.0505834101922909, -0.0952025766179358, -0.144213989856775, 
    0.0834979802606333, -0.137865110234016, -0.0806230072410678, 
    -0.124946411889084, -0.012684685245812, -0.327942126949755, 
    -0.0592088603965652, -0.198741620651214, -0.24363892695301, 
    0.184822327294265, -0.308511404915689, -0.0587815941751743, 
    0.0654889934026863, 0.0693891336400173, 0.0192631336681985, 
    0.0368525414236878, 0.225638280690914, 0.217367784489913, 
    0.079614899613305, 0.0896738110456581, -0.344378444071179, 
    0.280281537485424, 0.449898112846911, 0.215929963681856, 
    0.0650084137246787, -0.194468523685118, -0.122690267711856, 
    0.507802709511161, 0.414768508447146, 0.28022875903262, 0.41512607019739, 
    0.249911960244988, -0.300346614117385, 0.33332009993467, 
    0.605828919699398, -0.0361715881547732, -0.050716299031872, 
    -0.122587801850545, 0.566480838746979, 0.162097465488843, 
    0.0528276981658535, -0.146478424292147, -0.0425964942892576, 
    0.511566299422143, 0.151898267065545, -0.114679504926333, 
    0.107673196072047, 0.437806120826166, 0.0709962489029998, 
    -0.0271164361587789, -0.153402077893713, 0.190483864802448, 
    0.403229615116246, 0.010060799591071, -0.0799425141925112, 
    -0.127998153076457, 0.280087734173344, 0.156324516900211, 
    0.149013692117607, 0.320252760869132, -0.0605096453373216, 
    -0.33423619931899, 0.0479316126252511, -0.274516298127902, 
    -0.0167476284081015, -0.303024795742995, -0.0857952063405989, 
    -0.226381992488791, -0.202658920728816, 0.0457422410632145, 
    -0.105584899790674, 0.22200767499574, -0.07604113754172, 
    0.10407091479004, -0.265365467830019, -0.0279896523210838, 
    -0.108705831745685, -0.0599818889495944, -0.0872186109599184, 
    -0.0293706374270726, -0.205835562572411, -0.082643847877361, 
    0.0139478612886278, 0.107991531491548, 0.0886199486251871, 
    0.0428071834464834, -0.0194452376487402, -0.0208565526086155, 
    0.208340751850942, 0.199344138607564, 0.101973038789578, 
    0.184054727672423, -0.138037812102758, 0.543425610650776, 
    0.361346450555521, 0.0741870530172025, -0.137097720790564, 
    0.193894566621856, 0.603534734594535, -0.348249692410055, 
    -0.0452536815058599, -0.272842177609452, 0.313680087411995, 
    0.672779737172279, 0.266084613679303, -0.421806501049877, 
    0.0661892677405596, 0.0323719517792641, 0.517049705063183, 
    0.985790060537387, 0.189949619205405, -0.120943350090149, 
    -0.0543645197443542, 0.0243674230377841, -0.168739947823611, 
    -0.00694466743797061, 0.189144010404059, 0.197618137574677, 
    -0.399135547518741, -0.352523552454371, -0.048398187224989, 
    -0.160931214765502, -0.0968244845150412, -0.125178395731535, 
    -0.14481201152819, -0.0662874702216714, -0.141380798639022, 
    -0.0144735249291552, -0.0931634008107848, 0.155242304822645, 
    -0.145262877804749, 0.259153886623192, 0.161762838482793, 
    0.0659833370404624, -0.172292563985137, 0.167247252462785, 
    0.407753245368188, 0.223421277407198, 0.0565618501750607, 
    -0.130748706254857, -0.134376542324174, 0.51223004942348, 
    0.263136502117616, 0.0346040602121725, -0.0746272667671141, 
    0.357031328194648, 0.544119181062563, 0.437091802237513, 
    0.201070094274795, -0.167557343426996, 0.0836673899229487, 
    0.818001953494032, 0.255731723969583, -0.0529439577611691, 
    0.138463812513928, 0.566728512921792, 0.207260362937552, 
    -0.0503336482750189, 0.411183985053356, 0.472795544930216, 
    0.24014233147912, 0.137332587990643, -0.228542967215593, 
    0.214276536754957, 0.407983008151224, -0.0220268220969729, 
    0.176835400562075, 0.664628603384192, 0.251177994824266, 
    0.264992006087274, 0.330156539907187, -0.0845908942623182, 
    -0.0889593968935523, 0.0205814550595983, -0.0844504591062649, 
    0.290329542421869, 0.0328277439660764, -0.0864250629402483, 
    0.0502363074603733, 0.39868565955485, -0.0210851633318518, 
    -0.052392594804483, -0.103870483562618, 0.0408359450928082, 
    -0.10533245590198, 0.0181515114711156, -0.100106387453223, 
    0.0220796377613877, -0.0686335962990569, 0.0770726411008463, 
    -0.0411144192316285, 0.259829578752825, 0.0643631715776299, 
    -0.0183209104129039, 0.396989165522458, 0.27068029168513, 
    0.0717038170274807, -0.0354180562478455, 0.374598616258241, 
    0.239676540900182, 0.264535981368068, 0.428432431537999, 
    0.109152948932568, 0.185531248761867, 0.894263893488385, 
    0.203661759157558, 0.378015513210359, 0.793812101982923, 
    -0.334256401564231, 0.686458789894924, 0.640377510708859, 
    -0.300302261952054, -0.136528959122604, -0.126373124873147, 
    -0.12580384570369, -0.134212105057365, -0.0179312449824424, 
    -0.104147657211586, 0.126448259098517, -0.258446305938266, 
    0.120827260092521, -0.123667120567987, 0.18418167063778, 
    -0.0895119960180085, 0.0918248705824907, -0.282613620414751, 
    -0.0864768624161899, 0.0251090124406656, -0.0930347434518929, 
    0.174723003626999, -0.105969513376624, 0.0729142284196264, 
    0.0305903373532384, 0.0460111605975269, 0.0155607370982948, 
    0.0291537565660553, -0.00164524103856417, 0.0256271163361017, 
    0.0154974784516585, 0.0295459677078194, -0.0413364272592787, 
    0.0247830939595868, 0.0672898589843822, 0.0607144793491112, 
    0.0310299462187344, 0.0868665477371585, 0.088040102635614, 
    0.133099673405144, 0.130719211213996, -0.0217884970610758, 
    -0.280308794317507, 0.02530740505441, 0.684179643153924, 
    0.0927952651095486, 0.165524305687833, 0.329935396094278, 
    -0.182254589858487, 0.954588428556738, 0.0700134038280088, 
    -0.516152680796953, -0.160199270452753, -0.0422424157772962, 
    -0.156185181372131, 0.0899650622918683, -0.123435264782401, 
    -0.104224542861585, 0.0312725002957858, 0.417537360821553, 
    -0.0291875244544499, -0.0495751907434119, 0.0398603587378556, 
    0.082654473483406, -0.212184467786156, 0.160448469953855, 
    -0.191991177810661, 0.0537964187577259, -0.35820989104493, 
    0.0214398111165274, -0.401060038266028, -0.1777798363348, 
    -0.0685911421249291, -0.167662285432657, 0.219829796769651, 
    -0.0438311405089872, 0.0985776080912932, 0.297084414626527, 
    0.122391427948945, 0.0595798040615987, -0.105363996998835, 
    0.0784660605858354, -0.0134658580960379,
  -0.0984917784756411, 0.0462605825336433, -0.034877619532103, 
    -0.0141631462387682, 0.053706885734279, 0.0282454266542048, 
    -0.113699161247603, 0.202043897364922, 0.319209941672291, 
    -0.286602211284968, 0.486342467407557, 0.410154882920681, 
    -0.0911208546448004, 0.201099400208617, 0.221978416560106, 
    0.402731523680458, 0.989304394747841, 0.382495299644047, 
    -0.018710880736185, 0.0228182239428216, -0.251149998566419, 
    0.120158973703373, 0.163740602171263, 0.422146479267587, 
    0.446268555172434, 0.118023044578024, -0.01059659069824, 
    0.157315677449807, 0.225404408334407, 0.00460418160343951, 
    -0.0713562161176715, -0.0418292706499071, -0.0568064226072552, 
    -0.0519251093645312, -0.0441241143065716, -0.0532349270667028, 
    -0.0407089367492925, -0.0390604724537711, -0.0382080693303256, 
    -0.0172272503512958, 0.194006374876809, -0.0152566682743438, 
    0.24576888750393, 0.301091501644782, 0.13914815635466, 
    0.0697350404315037, -0.0614166062423388, 0.119747328661421, 
    0.470712371299037, 0.227227683271475, 0.198688569420589, 
    0.261559946615861, -0.00645794095622178, 0.729744297387952, 
    0.289315888025835, 0.0880900508669351, 0.122440669293748, 
    -0.292773934914673, 0.462394166116751, 0.46789425460633, 
    0.139204488537332, 0.116338421684346, -0.133416913264564, 
    0.142603266518632, -0.157204117165817, 0.0822743845593157, 
    -0.209578470693757, -0.0199596990335736, -0.329125307927346, 
    -0.187161266874965, 0.016921555667416, 0.0667695278987075, 
    0.158233866469021, 0.112662664599411, 0.147760142648321, 
    0.111991539473626, 0.143726662561182, 0.203100505028851, 
    0.12139526794655, 0.0369881206778777, 0.107879751961403, 
    0.169078459138912, 0.105522422504265, 0.114633340573386, 
    0.208809717523278, 0.146021650549857, 0.108573175321052, 
    0.192293738129544, 0.419856610041295, 0.435781886925299, 
    -0.233562731913316, 0.548080359991351, 0.482016388447943, 
    0.25869398260425, 0.274762433598604, -0.202409169695632, 
    0.82753761977698, 0.208887038389893, 0.00971610543436524, 
    -0.0173124919684596, 0.477949757399029, 0.254098747934234, 
    0.102832845989644, 0.116973643856881, 0.121404527017419, 
    0.0804302799665256, 0.230978437932044, 0.744547326815281, 
    -0.0918884037363137, -0.162358098292567, -0.0717802315257102, 
    -0.290573680268049, 0.000292271988794793, -0.407441494642568, 
    -0.159508996802359, -0.198660654573246, -0.198416720038343, 
    -0.187133421328892, -0.0472655497445943, -0.241600350856486, 
    0.141042776190119, -0.0327029978252962, 0.0448616545980652, 
    0.272279559719266, 0.242770716643594, 0.123814386616477, 
    0.036830218711595, 0.167606080058708, 0.172648322174205, 
    -0.0294290945462062, 0.344735528661246, 0.331981944096334, 
    -0.0494611958980478, 0.559743296095455, 0.642499099961529, 
    0.153399690984014, 0.0528342509320515, -0.315288899841303, 
    0.548551899260505, 0.660389626265481, 0.135096440056941, 
    0.269158593545337, -0.584477105593921, 0.431536834584806, 
    0.54721838175218, 0.40671059035911, 0.316566447376114, 
    -0.260740471021778, 0.875033411021249, 0.127654157342548, 
    -0.176748891524909, -0.0122625729990676, 0.141497344969436, 
    -0.0537917008429002, 0.0562239746104578, -0.412695634957763, 
    -0.128714047871604, 0.462225469124729, 0.353998540641072, 
    0.158270070868281, -0.22883665964515, 0.343257857245958, 
    -0.135121093292919, 0.0232122176345434, -0.39840621980499, 
    -0.075496021070184, -0.13448938016592, -0.196553392575082, 
    0.300057475859327, -0.327064156309187, 0.0861650616099745, 
    0.187287849556387, 0.0823758818224019, 0.114341905393666, 
    0.2591922078731, 0.217100202897386, 0.12135322172174, 0.153502564377099, 
    0.297753119580995, 0.291770657692047, 0.203282257715229, 
    0.184376388184433, 0.161741360737353, 0.119002720845826, 
    0.0829168162507173, 0.101012549916771, 0.114886645709034, 
    0.125620908785041, 0.149731238665377, 0.101009791470961, 
    0.0114167850683381, 0.0452432454674364, 0.0453571198010935, 
    0.0537782698041006, 0.0767083806688743, 0.0274421115473969, 
    -0.0253687161969996, 0.134915931922418, 0.0714431226866717, 
    -0.0275428124920835, -0.0755301038159316, 0.369915909116042, 
    0.174258221672564, -0.0730091788888326, 0.0118674027834058, 
    0.655668003808247, 0.142385352714092, -0.00813330485530514, 
    -0.0411997206798511, 0.570584875808484, 0.111352850541603, 
    0.0948507233941252, -0.451647725893378, 0.894023190455543, 
    0.430118967371005, 0.0941412274947313, -0.159752572211469, 
    -0.195520158329823, 0.32847445879752, 0.480738425724101, 
    0.31999049513543, 0.327216294173222, 0.353141984080285, 
    0.400405212924119, 0.355739415760571, 0.225959148074544, 
    0.214855773604232, 0.252662904652985, 0.0991261716797856, 
    0.0286298751502433, 0.467455015191933, 0.337198699775882, 
    0.143041240138969, -0.148207504948007, 0.280922094232641, 
    0.18173025738961, 0.131907503216904, 0.61681405010049, 0.395437656723244, 
    0.149973159443703, -0.210074364900623, 0.178191142405227, 
    0.187648333371223, 0.659106362025096, 0.435375000406427, 
    -0.0409268132903343, 0.0885899781236522, -0.224098580970684, 
    0.1320673240247, 0.47337307381453, -0.183368437348959, 
    -0.00355519096494233, -0.0541206894771989, -0.0502849979523345, 
    -0.0386129847649078, -0.050054878103407, -0.0190425483033147, 
    -0.0223008046137388, 0.0909921619439668, -0.137788411056117, 
    0.166427351260728, 0.197905092887087, 0.00185166217426848, 
    0.259576407239248, 0.276534856797393, 0.0930129843861539, 
    0.28032043398467, 0.358697595151384, 0.078844703732185, 
    0.0242973919324904, 0.199172587846141, -0.30615412819328, 
    0.532358054676283, 0.547770588873117, -0.0769621826992648, 
    -0.257660227296165, -0.178682743671264, 0.256890443096468, 
    0.584344307119009, 0.321329761588167, -0.10278917913036, 
    -0.196293271202978, -0.119942526197114, -0.19139493168954, 
    -0.0988393368417482, -0.220878669190116, -0.145088152814675, 
    -0.121106747356462, -0.128802483996521, -0.111586568252068, 
    -0.0070866500068222, -0.0317330814573044, 0.116328287117451, 
    -0.105328624794328, 0.107376837746423, -0.196587499602445, 
    0.00968365546077202, -0.062175246485008, 0.0517155757241617, 
    -0.224594150255178, -0.0240663971421609, 0.0381837781945421, 
    0.038537385642214, 0.0194809054755984, 0.0395877571179895, 
    -0.00596678688606704, 0.0139166968200884, 0.0194059101251623, 
    0.0185567238899909, -0.0156131501807651, 0.0372332784405574, 
    0.103783499786525, 0.169042358335553, 0.162002041326152, 
    0.117612159249609, 0.0652842267760193, 0.133052433429469, 
    0.366780895231856, 0.15696163198782, -0.172207629582566, 
    0.0946738387295605, 0.363011343509911, 0.335606656077765, 
    0.386177773090767, 0.276235145955459, -0.162413798617272, 
    0.778066442721222, 0.365510159042896, 0.00328308881707383, 
    0.310058904945683, 0.502191269672574, 0.0839287283959849, 
    -0.134352351736021, 0.322565013114409, 0.238870586662072, 
    -0.171800090218693, -0.251251450406652, 0.0543645128806907, 
    0.356104238874451, 0.000802935915491056, 0.0317368228263287, 
    -0.228954238307418, 0.256006710319215, -0.141422274152271, 
    0.219766554380853, -0.301830326670378, 0.128476579758939, 
    -0.522001726648828, -0.0739917746876908, -0.237968759619115, 
    -0.0752262689937881, -0.0343106919321253, 0.0995671576079357, 
    -0.0248134054225743, 0.203557241218755, 0.0393389344258208, 
    0.0613580025893055, -0.0779709551727148, -0.00498349620206287, 
    -0.1271372759526,
  0.153148688931448, 0.176806524799648, 0.135747317691477, 0.302705148592062, 
    0.231660665596582, 0.118888888758207, 0.338485685713905, 
    0.303978042487761, 0.23328602259534, 0.406225895614511, 
    0.242357856559938, 0.325849915912314, 0.769080526535381, 
    0.27669275028383, 0.142052860631095, 0.233038252335514, 
    -0.000773650045140545, 0.386011944587274, 0.209302879126036, 
    -0.196903649043576, -0.179748225081111, -0.1727172032673, 
    -0.146980814706119, -0.187426070172281, -0.106880564005055, 
    -0.212850066191394, -0.0365231308660068, -0.204293344404918, 
    0.0891424828786196, -0.229931054236686, 0.0612668907124442, 
    -0.0941526706953514, -0.102529658118046, 0.0424634590695836, 
    0.053908236068979, 0.103164715913775, -0.0754044194638529, 
    0.0448325572685401, -0.140980268574052, -0.0465594106634956, 
    -0.00220055061122933, 0.0603351358229268, 0.081020854474879, 
    0.0762694503409263, 0.0779433662793182, 0.0776120484369626, 
    0.0937288968725829, 0.10457128752918, 0.0708393949708779, 
    0.0961585869604543, 0.202324877879937, 0.0215269103886439, 
    0.112690785505269, 0.486644235894986, 0.175575982933351, 
    -0.13405345250715, 0.222738370653224, 0.453061417000232, 
    0.0631990505361594, 0.0509122206144093, -0.15785051637199, 
    -0.0571104884372547, 0.229635678344034, 0.769714398242929, 
    0.0149693704774313, -0.307371492239308, -0.00858476551288774, 
    0.631059041096109, -0.0592436179185864, -0.0134544450167817, 
    -0.187612366505011, -0.350987402637323, 0.00461889551527624, 
    -0.528094449171574, -0.296915697970426, 0.0975698173056008, 
    -0.327972526335551, 0.0684525412319393, -0.368876026278413, 
    -0.197243687585035, 0.0307739060137862, -0.055182524484672, 
    0.101884509796536, -0.0358350022279769, -0.0534793332809956, 
    -0.0120570708375325, -0.096298114654961, -0.0463209691651385, 
    0.172627932709087, -0.176939953016568, -0.00394775453978136, 
    -0.0634622198406097, -0.047750465632591, -0.0539252090662058, 
    -0.0510373851015201, -0.0616876438026303, -0.0337313785102607, 
    -0.0269628635126027, 0.0817208491139032, -0.15826108611808, 
    0.114462007566959, 0.199751268954946, -0.0651522442952655, 
    0.125820053518471, 0.342702957195907, 0.140546575106087, 
    0.0308156316888111, -0.0830059714459177, -0.241078823750197, 
    0.213896266753754, 0.531732158250789, 0.329224578463804, 
    0.119166621673196, 0.15172409776492, -0.271442611877118, 
    1.22921078620332, -0.311180438459862, -0.332336179887583, 
    -0.0484274417639647, 0.660395296965977, 0.105090258461593, 
    0.0870787535679913, -0.14532905099951, 0.152580565379904, 
    0.0398746806831711, 0.000160510883628104, 0.039295421956887, 
    -0.178706459930802, 0.062043721612364, 0.0792987528962321, 
    -0.0947626127488247, -0.0508175112336228, -0.13570501698383, 
    -0.0315227639084636, -0.118005331806316, -0.0636051887948722, 
    -0.0669460782910473, -0.114457613242613, 0.0571605577811548, 
    -0.145178375932843, 0.128305229981732, 0.091248433857408, 
    0.39213301085585, 0.23646896893533, 0.0428422151052316, 
    -0.230567132727725, 0.227184868312273, 0.44476266069009, 
    0.215898231211556, 0.0953502436067481, -0.0973117512296352, 
    0.348630904554934, 0.426580720345785, 0.120312463225111, 
    -0.190830726894954, 0.20577480627243, 0.765646423285353, 
    0.420067717171496, 0.149618735796829, -0.316601568217526, 
    0.47517885197395, 0.674691560362541, 0.168449731420989, 
    -0.31209814030662, 0.29185835404184, 0.474601768203178, 
    0.170886417716442, 0.0580223081678263, -0.153311845872624, 
    -0.0527127146456049, 0.319625793001607, -0.00766494062919308, 
    0.486161492122195, 0.331724775794528, -0.207807109000688, 
    -0.0281851920937928, -0.0578170039992419, 0.528644709673197, 
    -0.0450233006747818, 0.0158077183458251, -0.0113849845183748, 
    -0.244557625132797, 0.164971375282879, -0.0614173418613157, 
    0.100364715826834, -0.147733901815084, 0.0570187749787232, 
    -0.106830909533955, 0.0546176538664595, -0.312723665406779, 
    -0.00101863749167787, 0.0657465584513049, 0.124904707772637, 
    0.183573186075097, 0.239698677969202, 0.263993106081943, 
    0.238289062680007, 0.203872533901877, 0.227502908709124, 
    0.284509521574214, 0.286325053161664, 0.253162025880907, 
    0.241165070072686, 0.2453595929743, 0.236453706937572, 0.215298766742095, 
    0.178995093443802, 0.171539182631592, 0.258744557368656, 
    0.265606356341026, 0.149724200439105, 0.120686377436735, 
    0.118047528345575, 0.103021270249272, 0.0977043269060882, 
    0.0945320682448065, 0.0995722088738019, 0.123739141227132, 
    0.112866327219825, 0.0759110936282485, 0.115193177321906, 
    0.139835520409006, 0.172586283950801, 0.20346190877893, 
    0.205923363569407, 0.155576797198246, 0.12488250113396, 
    0.286693725936521, 0.290068158353365, 0.0761099180785784, 
    0.0145099626719668, -0.138731191719348, 0.666681982707218, 
    0.273455337921864, 0.153755241350294, 0.271589291848149, 
    0.488964589204259, 0.768223861957285, 0.20805953096705, 
    0.0491018912308004, -0.0425366505680964, -0.233576798495382, 
    0.11480517846985, -0.06583991514182, 0.0654594878135307, 
    -0.105873044672109, 0.0113541965480871, 0.0264033190218237, 
    0.0738401714066642, -0.228027175855502, 0.0329092803040243, 
    0.123041263361587, 0.163804678268592, 0.135640023923975, 
    0.253986342116312, 0.348240596165581, 0.217027448326061, 
    0.106908173816545, 0.229535264439747, 0.269389311293718, 
    0.070366868399798, 0.0810008490272712, 0.044971508790268, 
    0.0296992494799673, -0.122212105665164, 0.0409094629250106, 
    -0.0645983670266006, -0.0440726322389007, 0.020136541233179, 
    -0.102894591916873, -0.0981017529967718, 0.0697626594208107, 
    0.0905770763839521, 0.173334289602873, 0.132679093737126, 
    0.078734315221795, 0.274105586398113, 0.059053480299247, 
    -0.165574514358946, -0.22550853476568, -0.238966325353067, 
    -0.19879524260713, 0.830216797618145, 0.32722516858624, 
    -0.104421605818023, 0.0157818614564317, -0.464334235587283, 
    0.151584771025888, 0.16665666899927, 0.421989678596982, 
    0.958372494647963, 0.65376764692762, 0.184483138428164, 
    -0.309487543013358, 0.416729263645456, 0.413483644959071, 
    -0.0561972675447301, 0.0205912166119043, 0.838369569237018, 
    0.298064216776467, -0.00563754281297278, 0.0442610982878463, 
    0.389350552551808, 0.345141100487188, 0.128206790079475, 
    0.0541081232379711, 0.164848135031565, -0.14533107842498, 
    0.240123955114181, -0.113171449490432, 0.645597330639871, 
    0.619492010834095, -0.0714632810199075, -0.135953510467944, 
    -0.0172764197452493, 0.467946024564452, 0.110513828005222, 
    -0.0254637476967245, 0.605368067179002, 0.189305264611804, 
    -0.0458928948081649, -0.0997541899397698, 0.048892835697411, 
    -0.00694002624013559, -0.0248990040122556, 0.0405136751699754, 
    -0.0227104497415591, -0.0451337470441075, -0.012455868704584, 
    -0.0841021219473898, 0.00350155788628561, 0.0278457246492458, 
    0.257950168690574, 0.222750690599779, 0.0942120802928429, 
    0.104290353911316, 0.235186735563822, 0.160758903365656, 
    0.0972056947410679, 0.221200841849145, 0.247370324946816, 
    0.183824052362208, 0.142214683472581, 0.135837382622789, 
    0.139700484525608, 0.132457134931237, 0.123868398460814, 
    0.123265595830821, 0.131470946661929, 0.139900475865297, 
    0.135589296836911, 0.127057432351643, 0.103435391033658, 
    0.0962497318373174, 0.103367080601665, 0.106823554908524, 
    0.11309665684457, 0.146080458371303, 0.104244559957967, 0.0106355321336573,
  0.161859921490715, -0.342854341504977, 0.692735817579442, 
    0.583329211457404, 0.116906941496558, 0.765832298400191, 
    0.585968418586323, -0.392272815064802, -0.33613597223849, 
    0.129692677243962, 0.341121801467437, -0.00944288713748949, 
    -0.0573574520013672, 0.116630702622687, 0.287288559168522, 
    -0.136899756253741, 0.0495563663540869, 0.439381008337254, 
    0.186014835001801, -0.0383491685453256, -0.169933248323586, 
    -0.23643541368646, -0.00661827904092041, 0.0556710930699084, 
    0.253776113926995, -0.0766750585942732, 0.26093494448513, 
    -0.28449391085945, 0.107244385240063, -0.349549870579038, 
    -0.0736885021240264, 0.0564731722604249, 0.172981405897469, 
    0.170328292476732, 0.158232405366469, 0.157226027622448, 
    0.149329947087596, 0.137806988332372, 0.177801291711354, 
    0.204639087687167, 0.11001359433053, 0.0574418074245106, 
    0.0908606083471283, 0.116265374933356, 0.112149145408233, 
    0.0734339004565737, 0.0905829235839208, 0.103194612118075, 
    0.106937792067741, 0.0548661178507614, 0.0937618341357238, 
    0.0911362283043281, 0.0926601458599252, 0.201621454577083, 
    0.204997560365567, 0.104111752544834, 0.0146430813379572, 
    0.139663478600445, 0.338158508272709, 0.159398926095005, 
    0.044102597759213, 0.068501598174662, 0.582842370230984, 
    0.201412754846595, -0.328097137673441, 0.341965321739853, 
    0.673088062548724, 0.159562556904557, 0.00619587193859805, 
    -0.0740949223224874, -0.245005583323568, -0.0145489989802483, 
    0.684462799394669, 0.29813774635278, -0.0853208495845577, 
    0.415504992917157, 0.348485672515987, 0.0677285853763041, 
    0.138424270694648, 0.588008911704135, -0.0151316188837551, 
    -0.0526040663875634, 0.00699897576624492, -0.204405058732996, 
    0.0387774449668492, -0.041252194662605, -0.0732476003374276, 
    -0.0557165175525782, -0.0152695739074156, -0.0875025075696284, 
    -0.0995044032770093, 0.0107306933062801, -0.0546132166970744, 
    -0.101442767615316, -0.0594432800188074, -0.0154350191969188, 
    -0.0408778878016104, 0.0014821678337244, -0.112215557378697, 
    -0.0396538753076636, -0.0491808188887654, -0.081287790802977, 
    0.0804808616307315, -0.0976235224205714, 0.0711459024754575, 
    -0.209907580564807, -0.015079273862053, -0.0807339797349576, 
    0.0231572208029137, -0.195394046654174, -0.0263544724193525, 
    0.0562080711942939, 0.0666703516807274, 0.0452639214192309, 
    0.0339032635388392, 0.0493446016460183, 0.0969232405932689, 
    0.113003335664234, 0.0591106499088128, -0.0529848413857674, 
    0.0708809177679637, 0.304926591823452, 0.194870451359634, 
    0.017875379808598, -0.00906553014067588, 0.42421012131837, 
    0.407713177608857, 0.169007239143042, 0.00916653699859593, 
    -0.149304809346195, -0.284231015311616, 0.592603340720507, 
    0.482134808365695, 0.406420354129988, 0.255356660017805, 
    -0.102155836454131, -0.361235681376571, 0.764210986757493, 
    0.474017355082263, 0.181967009860518, 0.0541895121143382, 
    -0.114227002673651, 0.437417207852063, 0.682598614362232, 
    -0.228027975689847, -0.0150784827072926, 0.135635529686937, 
    -0.227551274795243, 0.469968212007461, 0.342860042234982, 
    -0.232392436394196, -0.185689757275684, -0.0897120122047558, 
    -0.198241210869586, -0.0154249289879826, -0.235185078372153, 
    -0.0547111663736753, -0.129873723897348, -0.0200127280362602, 
    -0.215060932920436, 0.142559437929265, 0.133431265894557, 
    0.0464320874631672, 0.0718878918639488, 0.144151183148551, 
    0.126074169118246, 0.283267707339637, 0.313436475047526, 
    0.146255885855095, 0.0576515463452655, 0.0122490906751618, 
    -0.0918544734665235, 0.0930001901401297, 0.300548218664472, 
    0.689960923286547, 0.384874017023099, -0.0789419183428268, 
    0.535801224648823, 0.411359101503134, -0.00336913765450255, 
    0.130854683505722, 0.639764783697961, 0.272364707906567, 
    0.117214956979649, -0.199352927077723, 0.0982106221148817, 
    0.295741081403832, 0.17410647699194, 0.841231686275762, 
    0.328930819700957, -0.139628544884069, -0.00125346994016239, 
    -0.110820472681573, -0.0345882268498052, 0.292990390713874, 
    -0.0276776638975833, -0.143028090708893, -0.0229496605748049, 
    0.21435732291713, -0.0799204971923725, -0.155211825354364, 
    -0.113994877863234, -0.152139686001186, -0.182126454830341, 
    -0.0987581096890928, -0.0631205455585893, -0.223610690327938, 
    0.0845230019388767, 0.0556067137725518, 0.133251874000372, 
    -0.372481970589992, 0.0238596759610524, -0.210694238266616, 
    -0.230252886652861, 0.0699891505871245, -0.130370044701032, 
    0.112582464275167, -0.154359102962983, 0.0910227059765509, 
    -0.347434909333454, -0.0741713031050384, -0.0202133785819552, 
    -0.0063630149117848, 0.0141872702592847, -0.00107667133322491, 
    -0.0152582432577471, -0.0306063401002726, 0.0243496945091203, 
    0.00900457160703968, -0.0243279619854652, 0.273442460307889, 
    0.122253646197421, -0.230034494619975, 0.28747411620887, 
    0.400110786910345, 0.161294521212544, 0.0733163973145167, 
    0.363916137600504, 0.30619860555461, 0.266183010182293, 
    -0.369430298274584, 0.734283842946007, 0.647167538765961, 
    0.316464075372423, 0.242854598877393, 0.908751747415087, 
    -0.0198197268860515, -0.132674735182218, -0.090968523695582, 
    0.651594511499583, 0.269854652525476, 0.040999401201192, 
    -0.111724375860468, -0.120596200209797, 0.322192241251482, 
    0.184910284976958, 0.103920667203379, -0.132084755249561, 
    0.228756296801166, 0.210822196167843, 0.0505891229822136, 
    0.195272295818967, 0.176824094654536, 0.0327793281600836, 
    0.0442315984758203, 0.218825980724236, 0.160432181911032, 
    0.115926613530575, 0.1123098813023, 0.0255193046934957, 
    -0.0283930975784042, -0.147055433185259, 0.120057385726911, 
    0.316023346101815, 0.138413157419116, -0.012755596822082, 
    0.015317555004632, 0.471150231827425, 0.106311190219082, 
    0.0040269533699541, -0.129259075984182, -0.0511037685370789, 
    -0.1016211551399, -0.0314681234373076, -0.0948639891277974, 
    0.0182092172197326, -0.120647506725945, 0.0236674756052266, 
    -0.137165287378492, -0.0383517913944388, -0.0258374979899113, 
    -0.0235597325440102, 0.0661458356343047, -0.0280809743454336, 
    0.00937313933799605, -0.0953104751994471, -0.0519841870584768, 
    -0.0150605279482399, -0.103682244205286, -0.0618533556113886, 
    0.032743274995946, 0.0548760234016387, 0.0811932597904951, 
    0.101739109455084, 0.0847235411474231, 0.0530721352560163, 
    0.0652757103742684, 0.270027592989613, 0.191338146369361, 
    -0.233942137108667, 0.240167281737639, 0.353238153506701, 
    0.119875474633863, 0.301360614913581, 0.254631071185612, 
    0.133049199644485, 0.747820202431599, 0.393203089461711, 
    0.00566963942078308, -0.198214452676398, 0.142617078213539, 
    0.301426551326315, -0.0807896400009987, -0.201656082806656, 
    0.0768581801018816, 0.343609183662565, 0.132259007402415, 
    0.117171656914291, -0.0912964386058354, -0.249499862496044, 
    -0.412788833905963, 0.085242407687105, -0.331931008728382, 
    0.0164043254970633, -0.372955660820749, -0.0749928412123091, 
    -0.189144055864352, -0.223759692535973, 0.186015460909175, 
    -0.33786394863708, 0.0596893959920322, 0.0754727276223416, 
    0.112476907669271, 0.0855646537333285, 0.113566337207088, 
    -0.00401231695512735, 0.0988394303679777, -0.0545907632788388, 
    0.0153482669122733, -0.0901633155193484, -0.0954771688177316, 
    0.0167847008918185, -0.0647210568082146, -0.0393372327776955, 
    -0.0151853442320693, 0.0159953463486489, -0.0346764008890862, 
    0.044063697050325, 0.249560819581429, -0.0930152092339273,
  0.422422697842266, 0.0462663789314664, -0.0888605264023776, 
    -0.129276588755862, 0.387175749042766, 0.383897464969548, 
    0.394903275357861, 0.497691617043445, 0.134322547529424, 
    -0.0449522220096332, -0.282815280942575, 0.517583105695104, 
    0.24087831790608, 0.332853563910795, 1.07136553819189, 0.20020368239136, 
    -0.346223086058921, 0.180395234243216, 0.870911408165952, 
    0.211354603559938, -0.213704144753366, 0.407441834129912, 
    0.52223735323326, 0.0262243752140361, -0.126571410889136, 
    0.045690419541656, 0.0184051582868612, 0.0943906609584978, 
    0.877084016446731, 0.129987235744966, -0.0696469477698121, 
    -0.107977641635662, 0.336714530562335, 0.0720706034782895, 
    -0.0585963823863237, -0.1222568840628, -0.186731961635876, 
    -0.0655222589515861, 0.375467300066931, -0.0800882742109664, 
    -0.229384025766575, -0.14883143279169, -0.18884378113455, 
    -0.103894426099077, -0.163270536691137, -0.130526715412526, 
    -0.0490527042021677, -0.144047449151719, 0.0210260800817591, 
    -0.165274289492123, 0.00462846683765197, 0.0784593180834909, 
    0.121752691323967, 0.0886235849604394, 0.0953553378159292, 
    0.103988509275745, 0.0953910039936896, 0.0960061025819454, 
    0.0942805517517632, 0.076233228099097, 0.0754752065764637, 
    0.0744877983860251, 0.0961892723867625, 0.0941630276014639, 
    0.100050672941378, 0.0806674744127211, 0.0804220910980009, 
    0.0837598365664182, 0.0979830711727007, 0.100620011386707, 
    0.0337021225189396, 0.00906875217370552, 0.0380614407166796, 
    0.00631427138889819, 0.0296753720987122, 0.0138946602134334, 
    0.0372325704391484, 0.033810373818177, 0.0383050669318032, 
    -0.0239520966347663, 0.0381465987380302, 0.0311439170115421, 
    0.0330819508882236, 0.0424858042184216, 0.0452680714418337, 
    0.0168755046716067, 0.0741999000941843, 0.0680488093612236, 
    0.122852350373452, -0.277384584299717, 0.73311373131451, 
    -0.0361673210247442, -0.391439667098734, -0.047482306008105, 
    0.271118744471728, 0.729277931363795, 0.49125470913594, 
    -0.313175913415334, 0.594862493477157, 0.774110569754429, 
    -0.0898144101949675, -0.051496936538914, -0.0793275433200188, 
    0.00454206352050947, -0.0351309571324103, -0.0476156764214577, 
    -0.0855183372884447, 0.0599922069782277, -0.0545884845381329, 
    0.107117200369561, -0.21141889069665, 0.0936482295248947, 
    -0.399959569382993, -0.114774641120875, -0.0782961269886131, 
    -0.0929671555298573, 0.0437516507731859, -0.0433570071192135, 
    0.0235263424844513, -0.406496823507699, -0.0385948507753675, 
    -0.284987743299053, -0.235705781312763, -0.133391980542815, 
    -0.257677960146101, -0.145946258483896, -0.16005719192768, 
    -0.179196202079463, 0.0880028659462233, 0.00522004894437142, 
    0.793600905797422, -0.590570428189695, 0.442604723397089, 
    0.493811262161847, -0.14421978374561, -0.0937138236404879, 
    0.0843170785394172, 0.0772083868994723, 0.863526340655433, 
    0.204823181630014, 0.072487640418831, 0.0607161930596579, 
    0.151552362456217, 0.236697570465338, 0.26133262355502, 
    0.208844703475824, 0.0825675864436551, 0.0430942086300695, 
    0.216999904877989, 0.171305752129012, 0.092280634907112, 
    0.0886474239637681, 0.0954259334326654, 0.110658682164315, 
    0.123464326012875, 0.0921037645176475, 0.0526894771287703, 
    0.0658388945897322, 0.126912478643574, 0.170431745836552, 
    0.184882469925465, 0.129925153161649, 0.160256735650984, 
    0.203846843502011, 0.126199485808902, 0.00510803871091059, 
    0.301658118709681, 0.214334812335572, -0.15017337131593, 
    0.0287516935976493, 0.579430423679102, 0.10028242104204, 
    0.413331015128509, 0.680433431748107, 0.047773826837268, 
    0.134863436493165, -0.447571382776602, 0.0308882092972625, 
    0.749481118392281, 0.233669505819348, -0.135403113692343, 
    0.179773176100911, 0.576962231016958, 0.291371768027321, 
    -0.245088662976065, 0.732494396758141, 0.352978243693492, 
    -0.0482858725949346, 0.392226663940484, 0.537176904188469, 
    0.103379238841841, 0.0817157698112626, -0.127869626632184, 
    0.156378386071768, 0.274177820799197, 0.119248588098222, 
    -0.00818962759719276, 0.122332882798817, 0.263335003217097, 
    0.116997361829488, -0.0880826454391569, 0.0656662886854921, 
    0.790565886545669, 0.020259193797632, -0.111955771773459, 
    -0.00457019330988513, 0.463205952613954, 0.365105170537876, 
    0.271892345138783, -0.194726827590383, 0.0188565533342579, 
    0.312852531328893, 0.515407223330895, 0.171774081238568, 
    -0.135927297707954, 0.0385353160150436, 0.325445444351357, 
    0.159492469388489, 0.664535695032802, 0.252137585234727, 
    -0.140238830757639, -0.0412516279832849, -0.0114760645810231, 
    -0.0434973651974602, -0.120876079077388, 0.0930373761171633, 
    0.0352300837271897, -0.0452077205403628, 0.0449848669419203, 
    0.0584443182768984, 0.0408516406788179, 0.0403427907678713, 
    0.03933002135387, 0.0250094080401859, 0.0238896320441563, 
    0.0728368199686159, 0.0830658802999765, 0.0459626164428192, 
    0.0389999155030895, 0.0796967404020339, 0.0136462028492101, 
    0.0288857216204132, 0.0408250883059652, 0.033128754309725, 
    -0.0738285917886892, 0.0298827846560377, -0.0772417690425529, 
    -0.0572886794515767, 0.034674977682394, -0.0602776719738551, 
    0.022836806202526, 0.0707297686822011, 0.11133301753838, 
    0.127189024936477, 0.111152776807255, 0.094568990000414, 
    0.147317084811913, 0.17777021635957, 0.0961868423322957, 
    -0.00403169235692109, 0.350471059163182, 0.247193403709872, 
    -0.0490252862201594, 0.294939433938699, 0.447556617695728, 
    0.157118046942692, 0.012179651593307, 0.349723098706967, 
    0.248309240703483, 0.224559131751023, 0.697073545273582, 
    0.327339905477165, -0.294051550705001, 0.298694219786273, 
    0.650545197800951, 0.497418474164933, 0.194309152351255, 
    -0.347670966015672, 0.0595967925618284, 0.427642635456834, 
    0.213368489775129, 0.361821263676374, 0.254670118707385, 
    0.0125874043003723, 0.380203469942731, 0.260850029377809, 
    -0.00683113895396174, 0.0373007694883904, 0.458419780286051, 
    0.0244269228656116, -0.0267627531847889, -0.0328476575103138, 
    0.0152819071746045, -0.00994481692836266, 0.00373172496065274, 
    -0.0120709632454363, -0.0514735651740835, 0.105299152892803, 
    0.0873665334619614, -0.0513910682640621, -0.244350894499842, 
    0.446666681390514, 0.244763770885124, 0.00739228128479848, 
    -0.116310588853942, 0.56383072928861, 0.383223834004112, 
    0.045914700051261, 0.804534813819094, 0.228579401340286, 
    -0.23152785826922, 0.478035905233794, 0.633847790080161, 
    0.109698552529131, -0.161198528355243, 0.340755824795038, 
    0.758422384389545, -0.0933786712096789, -0.246553742090373, 
    0.558136061549036, -0.00732056583372477, -0.112899797524202, 
    0.0430711343123851, 0.15932543668997, 0.168430861332031, 
    -0.24242353215713, 0.0111473919161899, 0.231653282631017, 
    -0.168152911621174, -0.138173286228006, -0.193832360518177, 
    -0.171073724364378, -0.054558143419595, -0.155721388019344, 
    0.0425736440749589, -0.144442465536824, -0.037930575177858, 
    0.11693844634133, -0.108550433282844, 0.110885107488862, 
    -0.049459385682109, 0.068759558999863, -0.00121608632978301, 
    0.0939781315515981, -0.164940311516086, 0.0263509578406107, 
    -0.263999264443651, -0.143059380266444, 0.0145216969246951, 
    -0.172244582059939, 0.00683835414529457, 0.023533256340009, 
    0.0122332320271088, 0.0995512213185708, 0.121219537503491, 
    0.0684122127685604, 0.092917049868477, 0.116117081832189, 
    -0.070346961802034, 0.163184167631409,
  -0.0555484077468518, -0.186727459126981, 0.0987155761989621, 
    -0.0556819460855163, 0.0753876900430405, -0.0609286898864894, 
    0.106568690888284, -0.043693055238797, 0.146961734250629, 
    -0.169939190584152, 0.134756327306012, 0.048646939190167, 
    0.0201454542873268, 0.339033368186952, 0.20928059963521, 
    -0.0164761795344077, 0.0668249256906807, 0.54167751651547, 
    0.15162762616315, -0.447193952560117, 0.222834647553772, 
    0.769707246684049, -0.0124835807516848, -0.260135372990092, 
    -0.120532489632038, 0.672078013329601, 0.208368929016709, 
    0.0678686764049411, -0.0465082558357485, 0.027541200917096, 
    0.0170473081964057, 0.766716903759318, 0.32035483951403, 
    -0.00487188046711387, 0.495446227388427, 0.24411803751875, 
    -0.107103740831468, -0.0225649608702098, 0.562494657523175, 
    0.0934290343446343, -0.0181407570171984, -0.17577199550779, 
    0.0920024004193953, -0.0581195804599224, -0.111238296735987, 
    -0.11176548893649, -0.0920978635006834, -0.0971405394286195, 
    -0.34753465446318, -0.0352129517882355, -0.249041680857575, 
    -0.165694792262982, -0.161310220635934, -0.011791224452691, 
    -0.156343813887165, 0.130901331225262, -0.283163284169793, 
    -0.00430224635850804, -0.212172221663116, -0.168623214320942, 
    -0.00405350823364102, 0.0476989659045908, 0.103076834023035, 
    0.15335154958201, 0.146184556692616, 0.126836499093877, 0.14018252417256, 
    0.16079362071116, 0.15037693517624, 0.142989017333913, 0.174920875538983, 
    0.181680946257808, 0.181051915304341, 0.184987297751813, 
    0.175406387281761, 0.15439567824559, 0.170453253802018, 
    0.229478617619106, 0.173283358945229, 0.0593460008000348, 
    0.0752558622650606, 0.318104233464134, 0.275282197181321, 
    0.109241995908983, -0.0818752770982289, 0.236698413380437, 
    0.452422990126404, 0.180065681431615, 0.0663293591666891, 
    0.0627026629665574, -0.057465778410838, -0.138218319201467, 
    0.80245377403673, 0.253280865651342, 0.0170408075321391, 
    0.341847428297672, 0.581583088429807, -0.368520587777223, 
    -0.484450230411464, 0.158648952710854, 0.335073952825387, 
    -0.150118918267272, -6.74046659596139e-05, -0.0698714945610482, 
    -0.00442967637418749, -0.21973465336661, 0.399692927479846, 
    0.166495255287464, -0.324964283922258, -0.0654852453826874, 
    -0.335785770190722, 0.106459910900607, -0.286240258312545, 
    0.0878785766160887, -0.219136788518318, 0.114446325400508, 
    -0.37050533495756, -0.0177183889770072, -0.327744478718185, 
    -0.217497272330425, -0.0445689302394342, 0.0986904675537526, 
    0.0218935525388694, 0.0587930319277099, 0.0114406501357557, 
    -0.0156747496357579, 0.0610699640512387, 0.0678196077664414, 
    0.090246681416785, 0.0078708889304907, 0.163903107720873, 
    0.132951990560964, 0.00731119914296696, 0.198599000347343, 
    0.371236256869575, 0.169528631968364, -0.0321097105332408, 
    0.282875526957838, 0.403735458061439, 0.160714473188434, 
    -0.291668637889985, 0.279915002480148, 0.485728374626899, 
    0.0457812039210295, 0.0857758583201383, -0.323119560836613, 
    0.290609315913012, 0.512524919007856, 0.201974162588742, 
    -0.132986209364903, -0.0250010618829302, 0.336901887451989, 
    0.353347730529744, 0.112252776264784, -0.205557999339143, 
    -0.0236630288321575, 0.327820065956947, 0.14987544355371, 
    0.209889219518213, 0.524187730383437, 0.117977367692893, 
    -0.00272895718888688, -0.0665388819597842, -0.0325929125838898, 
    -0.184698248031225, 0.0325883705159394, 0.0460897676170125, 
    -0.181440693323631, -0.050375803148363, -0.0773142411189115, 
    0.0424360528279202, -0.122402052592786, 0.0917006385645227, 
    -0.0780376632721422, 0.0703092269611377, -0.0188265209851607, 
    0.11459271136959, -0.0771766213044859, 0.103583574101039, 
    -0.212217941146208, 0.00919283696299528, 0.00402048906269661, 
    -0.00405443035108946, 0.0127753491374867, 0.0463755834235036, 
    0.0603901061305742, -0.021682090835916, 0.0535554295621412, 
    -0.030575152537117, -0.0346578484186069, 0.0774839397130875, 
    0.0584080709554158, 0.0591121497515258, 0.167122736763933, 
    0.128716285982374, 0.0545583152020561, 0.132064277114099, 
    0.163806023346524, 0.129807403397552, 0.0757486443777593, 
    0.103234159910303, -0.305230130646856, 0.316712629730584, 
    0.42766683390133, 0.269030441858366, 0.375729194467005, 
    0.312107285793184, -0.440346731299883, 0.261965080868063, 
    0.432676690790796, -0.0277868992833529, -0.0715151275085759, 
    0.151294469520488, 0.12530062831816, -0.227710824849529, 
    -0.200763023256998, 0.121208468213048, -0.161737168711812, 
    -0.159832458614791, -0.0677153855601466, 0.0570755782125721, 
    -0.349774341415308, 0.131848666664712, -0.195678532845947, 
    -0.0205897521986403, -0.251534856679933, -0.0928254670587083, 
    -0.140224105421578, -0.015625741115162, -0.366280729381597, 
    -0.0108650550149887, 0.0454581069284965, 0.112553453241753, 
    0.158122846448909, 0.142965263950145, 0.0983984458802671, 
    0.115109620545891, 0.145812782376891, 0.0982818208242056, 
    0.0346804198536957, 0.0641515850445893, 0.0257890391925669, 
    0.0543966504533351, 0.0172114866178195, 0.0347266770105149, 
    0.102097652958795, 0.18762943027503, -0.0470458098046789, 
    0.240588106705673, 0.189225833170369, -0.0663395912384258, 
    0.404121700737947, 0.38385243212292, 0.0895651273173902, 
    -0.256388315225457, 0.524186015759995, 0.342281515930817, 
    -0.21017265441082, -0.221394880044259, 0.597000654868991, 
    0.393904447478997, 0.184805296784601, -0.080607147609458, 
    0.258642882115393, 0.330865300358817, 0.0819417747961467, 
    0.266350928257259, 0.500417419344192, 0.292905447798111, 
    0.184984459990163, 0.32184932928668, 0.435144961582473, 
    0.346844324568777, 0.239784716112325, 0.131892941498601, 
    0.0422791843747667, 0.0978666671002943, 0.281443919263882, 
    0.0955575518799246, -0.320505340183624, 0.145128879452451, 
    0.555560817768571, -0.0458343746976108, 0.143389823775083, 
    -0.480441758683193, 0.305432429030445, 0.531417116887995, 
    0.270583731185973, -0.032107704980044, 0.278836961017861, 
    0.23244640807389, 0.0953697455129369, 0.676304838555675, 
    0.405494446986718, 0.170916116291385, 0.274253869909677, 
    -0.29113485785981, 0.500856472230112, 0.585728648186925, 
    -0.202053421787339, -0.205079135800705, -0.0158306209472698, 
    -0.0934592103484277, -0.0625494568752208, -0.0846097613485277, 
    -0.0358698571023515, -0.0938789674640188, -0.00709285164377355, 
    -0.0679316062168268, 0.0612796368186357, -0.055135340610893, 
    -0.0341086274353752, 0.565716250149506, 0.12101271486219, 
    -0.0274225573566472, -0.185895950039351, 0.529584654633596, 
    0.25559211076776, -0.14488517846217, 0.232345103060543, 
    0.632033143073393, 0.243754154585084, -0.206836078685914, 
    0.397570379032088, 0.510367613693394, 0.149867261108697, 
    0.0288136344272734, -0.210960646961028, 0.334023643303379, 
    0.547746779957084, 0.250616693602265, 0.168548793305227, 
    0.202218977668422, 0.290621030466304, 0.301109753675583, 
    0.195408293537662, 0.111792788578098, 0.183505452811514, 
    0.272636986231631, 0.129110071505349, -0.143125067296577, 
    0.283375049620964, 0.409125323010402, -0.0787864468294046, 
    0.0117638997102502, -0.155411150003552, 0.431515726070571, 
    0.173881267459646, 0.123651918362103, 0.136183208153518, 
    0.0800837263182203, -0.139466292842195, 0.0364700107494795, 
    0.361340986138315, 0.357443576141048, 0.172256896632706, 
    -0.0983952795219905, 0.270902431209358, 0.27315978140722, 
    0.0605193764163193,
  0.0922726726802104, 0.00838822291320905, 0.170805105460149, 
    -0.176454064329803, 0.114835905717333, -0.202263076800259, 
    0.00586847775880264, -0.0972768705525803, 0.0665854596200316, 
    -0.171084755737134, 0.000820722972086033, 0.0283097064702166, 
    0.0346359218269456, 0.0245962875687716, 0.035076971380477, 
    0.0292246322020105, 0.034477457249238, 0.0340955599835364, 
    0.0352333321455167, -0.0482734815915542, 0.272631222681481, 
    0.188687588825683, -0.0303274051511207, 0.322904761369298, 
    0.336403760405651, 0.132272995916405, 0.0361545991360835, 
    0.173160154826279, 0.273734006823646, 0.333907348075495, 
    0.162169768449218, 0.231505645713979, 0.790252492282688, 
    0.321517437826871, 0.0910662751593271, -0.0176075742440841, 
    0.63162412177661, 0.216401592078392, -0.158581576992714, 
    0.323710294215936, 0.445603314161934, 0.200716647707919, 
    0.105565436155651, 0.0894358790985794, 0.0878089899652059, 
    0.072882708621192, 0.0728852031902308, 0.118356562967787, 
    0.0910062928912419, -0.00427226346528284, 0.0931816247730977, 
    0.262267132189222, 0.150864984451312, -0.0203683605049619, 
    0.178198247078076, 0.351118471587565, 0.285537138897786, 
    0.120152496327451, -0.16633550587935, 0.0375980656276646, 
    0.292216012540058, 0.286395053144568, 0.602977860148163, 
    0.293605762005389, -0.146057879770366, 0.0285920606421406, 
    0.766123665810065, 0.224068499992768, 0.0829454112978262, 
    0.280337027666436, 0.00993995610414143, 0.212964788435148, 
    0.486761550856944, 0.13896018609649, 0.0656898433463865, 
    0.129510120064925, -0.0592408831019376, 0.244879232215967, 
    0.135679258385187, -0.0356287088498304, -0.0926063208466725, 
    -0.258640770866052, 0.025744375753269, -0.101155612102205, 
    -0.00873105471649425, -0.129395640780498, 0.00685942243077964, 
    -0.137191122971317, -0.00307001699491405, -0.254282545362549, 
    -0.0448549079023917, 0.038494543098812, 0.127353310350086, 
    0.1531054372284, 0.121605104325346, 0.0830654234288178, 
    0.172934153166184, 0.277742810932516, 0.141084233136736, 
    -0.0346411448164221, 0.121311723900973, 0.438471156374048, 
    0.215326250619108, -0.0177290246577958, -0.00825257944951069, 
    0.530449098040941, 0.476203147046741, 0.0814264977762926, 
    -0.12854945499131, -0.122781255062774, 0.601745898219654, 
    0.226867781633133, 0.0575015121821377, -0.10114747989618, 
    -0.131140805675615, 0.641682156813784, 0.0811924788091458, 
    -0.169013935294901, 0.133278112748638, 0.460034632773784, 
    -0.0812818357599519, -0.0537571733061138, -0.133657915336253, 
    -0.052399012086154, -0.0384458252514664, 0.00489337800049164, 
    0.0321514673844237, -0.0151320960586531, 0.0298733361880441, 
    0.00330804402184191, -0.0378126872760604, 0.0764403549023798, 
    -0.103052874194002, 0.00515903874019417, -0.0473705918608811, 
    -0.0162308873944922, -0.294396457221371, -0.0336547035816856, 
    -0.213405837762341, -0.241104388028447, 0.00121148632958737, 
    0.029109985540625, 0.0332413097899707, 0.0515378924738723, 
    0.0661839076821527, 0.0391294597961435, 0.0275240667449548, 
    0.0976875052999076, 0.0582935935314684, -0.00463415359250963, 
    -0.0148670210663878, 0.099271406297529, 0.163376040729149, 
    0.295564515236841, 0.468754761381237, 0.191999350563505, 
    -0.143864605945558, 0.104059829687134, 0.509206163383031, 
    0.268006821198612, 0.117942132799742, -0.19551644332426, 
    -0.0152904698463842, 0.738195925248484, 0.0560204906380337, 
    -0.0847584991025168, 0.056054346934955, 0.453881797426494, 
    0.765801910552361, -0.197518692207921, -0.271796637748212, 
    -0.0570746128804221, -0.169813672830708, -0.0387967418709863, 
    -0.193161942659055, -0.112927763899528, -0.152851592627465, 
    -0.25373193111257, -0.112838370928972, -0.184101254659293, 
    -0.00563791895896284, -0.087264740562585, 0.0757053191307937, 
    -0.0433754809563232, 0.127130107863539, -0.0356048202897027, 
    0.0817876861629268, 0.0051530754187403, 0.0903808953414656, 
    -0.0679998461284504, 0.0580802887864021, 0.0123888141271439, 
    0.0277428581674788, 0.0245903036150875, 0.037425207110943, 
    0.0137081023179427, 0.0370910608933151, 0.0320777099338349, 
    0.0543242888636623, -0.0410472486972732, 0.0779917013867525, 
    0.151498339160275, 0.0902513753557706, 0.0588491455264229, 
    0.185911112960922, 0.194000302820729, 0.0970841853160962, 
    0.394303329465987, 0.252247119531071, -0.212375314273625, 
    0.0994008907287891, 0.507975696975349, 0.10116872111567, 
    0.522352758326369, 0.796126145178858, 0.0685585136548681, 
    -0.060334379904347, 0.487343157663132, 0.0495943748142374, 
    -0.0411854240690379, -0.287672690901055, -0.0364017009199759, 
    -0.230964710112429, -0.196589319841763, -0.0284284071690883, 
    -0.0692043107274442, -0.105988326860732, -0.0594057334840378, 
    0.0432709819933226, 0.0167988184690183, -0.226052093962964, 
    -0.0267243018215993, 0.0621319255205556, 0.104596819000738, 
    -0.232504117807292, 0.116195823592337, -0.331687740469302, 
    -0.188662684511998, -0.0510449585570273, -0.342527875505514, 
    -0.0764158743305338, -0.00742690774957219, 0.0208318315414868, 
    0.00374438179920894, 0.00515940179256912, 0.0397006915512439, 
    0.055044104028034, 0.120434514618984, 0.154202379438403, 
    -0.222378263593869, 0.308897288922056, 0.295680739670638, 
    0.0473526007225545, -0.163173485790687, -0.0491882710474324, 
    0.496656839484475, 0.418512663905795, 0.14266402809351, 
    0.120107823879226, -0.125119517143586, 0.808111536835142, 
    0.0566389329928026, -0.0968609503568418, 0.00580526111993397, 
    0.301589792951438, 0.810375753623162, 0.436260178837, -0.325652047004123, 
    0.165509840282388, 0.567117216952314, 0.101229590820328, 
    0.0276790912977069, 0.219316632818256, 0.187135070256083, 
    -0.0398141593089973, 0.258721769746321, 0.460787721975255, 
    0.166155054777088, 0.0538240150373131, -0.151037334002866, 
    0.13530961529388, 0.229974177091427, 0.213519387466677, 
    0.514825685013189, 0.247007884756799, -0.0497239483735747, 
    -0.10769316754129, 0.208313162846448, 0.397576833519266, 
    0.44338082810696, 0.253615243514061, -0.115540168482421, 
    0.358948735886836, 0.578437658854196, 0.305921682668881, 
    0.256958353621888, 0.347440270716943, 0.126227372979228, 
    0.811529644164807, 0.181141605790399, -0.241227910650646, 
    -0.106120969235258, -0.00769435726192738, -0.141122115744756, 
    0.00327927581338196, -0.0752343531939077, -0.0914918733486381, 
    -0.124127572722341, -0.0889623842941264, -0.0833235063267485, 
    -0.188945784581059, -0.0079344219083199, -0.120440260859228, 
    -0.113112391817804, -0.00767304805786564, -0.115145410036158, 
    0.0256570662514638, -0.0703998585392964, 0.079987573648878, 
    -0.0693096881276508, 0.0740821047484248, -0.0109773207141827, 
    0.0260036758618536, -0.0168548076023062, 0.00920774957038952, 
    -0.00152427954587592, 0.00814594141865703, 0.0378605634034383, 
    0.0194491439067126, -0.0184688312703361, 0.0449427969647005, 
    -0.0349598673619001, 0.0569306497648832, 0.397740204888374, 
    0.161370796361683, -0.0406858635404335, 0.0989974473789336, 
    0.357444407598674, 0.144088045547887, -0.346320921657796, 
    0.351107150755749, 0.998652305043656, -0.11442800587643, 
    -0.0182574623451241, -0.233684975659749, -0.211871636485662, 
    1.10940709448145, 0.277771158545928, -0.151384632124532, 
    0.211408879123898, 0.310320975914659, -0.0387604845425199, 
    -0.0433658164553377, -0.0756757827117982, 0.126716752903409, 
    -0.368900346439427, -0.0565201234735206, -0.25067914598203, 
    -0.0993236548334676, -0.296940726788229,
  -0.0368951257787292, 0.0548945211195889, 0.0592176846393476, 
    0.137358878119863, 0.17884558152237, 0.0895393426174105, 
    0.106172742801245, 0.291272321394586, 0.136587117500654, 
    -0.00981051989281279, 0.108235544703787, 0.357541352092106, 
    0.064687841414376, 0.0569494120757615, 0.820586071419066, 
    0.342971772858863, 0.07894409011683, 0.0493004364492893, 
    -0.0650091383381881, 0.17186129365922, 0.583495505099672, 
    0.409705228724286, 0.705374126496176, 0.659762024352049, 
    -0.0878378549521486, -0.123236873364759, -0.498188319065153, 
    -0.286356746623394, 0.860173689845278, 0.674814958053372, 
    0.216828845750918, 0.0652899568373048, -0.098333579422893, 
    -0.0830882789514322, 0.239085569314453, -0.162610052310537, 
    -0.112868189882706, -0.0365569373394911, 0.00543030083141294, 
    -0.142264589256429, -0.16792103862202, -0.0384758631885805, 
    -0.277572049504326, -0.140435258652056, 0.0850041403502183, 
    -0.183703925380772, 0.10491340678086, -0.0509741787189883, 
    0.124188739190114, -0.0924344143883171, 0.25041433517828, 
    0.0891926582455524, 0.0413758173367706, -0.0816305174268804, 
    0.330245501661264, 0.11577021811715, 0.0173287539531888, 
    0.0356887736884569, 0.0125971643654922, 0.243820975694631, 
    -0.167344812572433, 0.262888228225793, 1.04941939784613, 
    0.175592945502474, -0.135023059031732, 0.423235793809864, 
    0.749939797096513, -0.110332277538907, 0.537833824323268, 
    0.33206983261372, -0.40500131530292, -0.117035213443508, 
    -0.130713316476973, -0.0997186701591323, -0.137634006209606, 
    -0.135182126331852, -0.0418608343337135, -0.129986178650466, 
    -0.121654877779223, -0.106847564839827, -0.0749573082270012, 
    -0.0377907332524512, -0.0354217367019362, -0.0472859965224821, 
    -0.0279114707598446, -0.042497356186839, 0.00119458737052339, 
    -0.0350815444793231, 0.0533546107461574, -0.0687398117636738, 
    0.0219953175913359, 0.0659811241763478, 0.0836973981260543, 
    0.0969394461135218, 0.109416532988926, 0.109236183980191, 
    0.107823789026933, 0.0998431986267801, 0.0703260700039285, 
    -0.140470577797444, 0.241608678951037, 0.442642237817459, 
    0.145694787183293, -0.108373309268212, -0.0960710585334514, 
    0.336857583727382, 0.580329714501399, 0.152998393778475, 
    -0.130179322552603, 0.012631312975792, 0.471864677601918, 
    0.133347587697269, -0.225137015415883, 0.306614252387727, 
    0.737800371283733, -0.00571535944990791, -0.391550794191897, 
    -0.0381398138729187, 0.625752352359933, 0.0868877209144514, 
    -0.165669844792332, -0.098680630930738, -0.458709602487222, 
    -0.186265844487054, 0.0432025982061366, -0.341270842281063, 
    0.0608051884226409, -0.0791702055942753, 0.0617512052256121, 
    -0.303826379501841, 0.0169181928663579, 0.104731723399, 
    0.103525101184479, 0.192085195510947, 0.224581005516295, 
    0.167125183760798, 0.161355000974243, 0.222155365318064, 
    0.200120691043678, 0.127781945719362, 0.149265724030044, 
    0.220480499367508, 0.17832752878639, 0.145769334976023, 
    0.321314949321068, 0.326409169683671, 0.147496852053444, 
    -0.0222821491419083, 0.376481438185932, 0.342360221967692, 
    0.14248179064252, 0.0976634057957841, 0.520108724536955, 
    0.208249123761744, 0.019045883985674, 0.901927811217335, 
    0.214660062154904, -0.11094453244619, 0.520885969213961, 
    0.272511068007941, -0.271760041364114, -0.0759774299617968, 
    -0.133844190095458, -0.132058594063388, -0.0416736781649487, 
    -0.0960801869389903, -0.114400795284781, 0.00589570278505744, 
    -0.203117066939795, 0.0508462041459371, -0.244255912740183, 
    -0.115747242247315, 0.0737241603848254, -0.164432196283473, 
    0.0926204011536285, -0.0995070956893515, 0.00474810936140474, 
    -0.0357634550470335, 0.0402210172252626, -0.159112267252708, 
    -0.00172205387089247, 0.0636295774357551, 0.0730355503738078, 
    0.0986345237716249, 0.105672659468263, 0.0824693892252389, 
    0.0891120373357169, 0.129339779480692, 0.0960103779195102, 
    0.0269939680978314, 0.14958289180643, 0.199774117279099, 
    0.120071432830576, 0.199860394165127, 0.382336820236122, 
    0.202950869018308, -0.0193348354481899, 0.277850506323522, 
    0.477006473291577, 0.241261125521196, 0.116451821888003, 
    -0.279505963420728, 0.174981125896337, 0.692057363455407, 
    -0.241648807582041, -0.310826865239524, 0.0116873058195669, 
    0.589546753415382, 0.0482241473163675, 0.189323020726687, 
    0.158193984512389, -0.520798740832224, 0.266982951363963, 
    0.218565428794884, -0.0915726312220029, -0.0520495273119634, 
    -0.0935848512334311, 0.352937648790414, 0.0381899187352787, 
    0.0089491832983279, -0.292075777282478, 0.00634950900521983, 
    -0.22807135782389, 0.00863777206804568, -0.225665480905884, 
    0.0131971834818054, -0.245517632473134, -0.0993908302865812, 
    0.0135527986184515, -0.208928830270527, 0.27345058051957, 
    0.0562067681379202, -0.135841678588289, 0.166320517033, 
    0.451435559123656, 0.134669381662555, -0.00356825158914872, 
    0.0046506668491883, -0.0516533030498054, 0.131008373732193, 
    0.432490201152903, 0.554895358085604, 0.309160910662912, 
    -0.115425778365898, 0.616801934695461, 0.358901090418049, 
    -0.230858587423906, 0.370179321680201, 0.575544977317933, 
    0.0228554918611778, -0.11397381693245, 0.0265517707819261, 
    -0.216207583652055, -0.0500077502692187, -0.11120025783444, 
    -0.13246330553125, -0.00588776817849726, -0.131931895653434, 
    0.0149395394647708, -0.130587004288999, 0.00686666833988615, 
    0.0826510837704493, 0.127806568171499, 0.173580721067817, 
    0.202360875663696, 0.151575726159198, 0.106490712788351, 
    0.217964047048487, 0.279859178010564, 0.254678027250704, 
    0.187339957291166, -0.147583452433209, 0.161949122004789, 
    0.52905934748659, 0.224024850035109, 0.0885965414603013, 
    0.159672743184927, -0.0942347690601327, 0.243843247631254, 
    0.772930344163609, 0.118140775876401, 0.0322745363387669, 
    -0.0967395969458661, 0.736875286296487, 0.0766460429719612, 
    0.0513615317346186, -0.207446706789033, -0.0414475692114558, 
    0.507309172392366, 0.370909444949461, 0.0437731784771695, 
    -0.0492877194905067, -0.18663104759234, -0.100517425276787, 
    -0.202495868574028, -0.0914917390748444, -0.108376990555956, 
    -0.126355033717617, -0.134664066181663, 0.0141250196869906, 
    -0.0677130008281142, 0.0184494875253275, -0.00286808331183033, 
    0.00206833281514106, -0.190462173064468, 0.000830477400887736, 
    -0.0596838640587566, -0.0961044474357826, 0.129908328873232, 
    -0.175218207977102, -0.0290169865216423, 0.0533582512669326, 
    0.0715484016919497, 0.0760253641791632, 0.079232840780496, 
    0.0813587653584006, 0.0999828901983641, 0.108922435785085, 
    0.064388111378796, -0.0141768040622481, 0.165568072019115, 
    0.186073616479505, 0.0600040031247023, 0.213822065409862, 
    0.353994179156058, 0.187532126834278, 0.139091150740626, 
    0.246247629199419, 0.136208103484638, 0.453735780933703, 
    0.452607014940783, 0.0228474607298232, -0.0040720150766535, 
    -0.153585298553525, 0.506861053421616, 0.318188416444762, 
    0.253892638406783, -0.0370521518271898, 0.445468361285572, 
    0.298410244519408, 0.000438474844882145, -0.0316924263097516, 
    0.117124012472594, -0.0714409995220371, -0.126819839234396, 
    -0.165656915996713, 0.021019411509811, 0.0935332310463573, 
    -0.119550193273131, -0.0441146546622149, -0.0118417384553663, 
    -0.238778740683115, 0.125824010491649, -0.105146091724611, 
    0.0455595222093555, -0.236772281695552, 0.0182475668603384, 
    -0.153986567313548, 0.017291888004557, -0.258752508655902,
  -0.108206292501023, -0.173146804660634, -0.0570528560170733, 
    -0.0985787071586817, 0.147860229183637, 0.0462203171376151, 
    0.0841624628033347, 0.252706325233699, -0.0494875865086646, 
    -0.0499496874805157, -0.0354007754776045, -0.127821023138633, 
    0.0594717384136444, -0.103512808903392, 0.0107838860720764, 
    -0.0740968314955199, 0.011921774187107, 0.0481881423905115, 
    0.190382789098482, -0.18565385656012, 0.0580757080554271, 0.333372907558, 
    0.234791879793241, 0.197447408430772, 0.288228265176428, 
    0.146300812625028, 0.000110146594891697, -0.375939071969131, 
    -0.105127660780973, 0.474299875188575, 0.392975787789537, 
    0.413634948954618, 0.501830388577189, 0.299800031712598, 
    1.03255030173385, 0.116562987807422, -0.257155364899361, 
    0.348730571694735, -0.0928054063456431, 0.763636552362687, 
    0.00138943010399917, -0.0602505505800152, -0.041584767840529, 
    -0.12972292274356, 0.14155813369708, -0.0251431197561221, 
    0.0188527317710904, -0.0638885982575651, 0.114811892592965, 
    -0.00934804284483017, 0.034295765730339, -0.0942352032084588, 
    0.0397593488654374, 0.166607998775486, 0.0603542743531901, 
    0.0347591670588273, 0.0372774492882191, -0.0689341519974156, 
    -0.0796680092546447, -0.0241230569320749, -0.197048066854689, 
    -0.121137849342895, -0.0700972145945511, -0.0382791509982491, 
    -0.104565711290554, 0.0773746744028736, -0.169774037026312, 
    -0.0365212842788231, -0.122296743118715, -0.163091388267658, 
    0.0265123127201458, 0.0644972254333656, 0.0570218758408546, 
    0.0930194094588376, 0.108731264212993, 0.0820400991990047, 
    0.0838513608556297, 0.128777917679729, 0.0967203494318962, 
    -0.0346861924729919, 0.162759821510894, 0.310057804734997, 
    0.151163134856795, -0.0384313763574441, 0.12962338897813, 
    0.415566155314257, 0.390463486519045, 0.152500570176592, 
    -0.245422364479985, 0.110180095866858, 0.578023084955686, 
    0.0975124322983196, -0.244740848873514, -0.0290606395275173, 
    0.529012655664805, 0.519630850045538, 0.516896764361001, 
    0.388961869244979, 0.00639491141860715, 0.7500419282045, 
    0.37242974188363, -0.222200885818729, -0.13865725434853, 
    -0.227327083011652, 0.643274791805986, 0.0057068250445626, 
    -0.0405152404953973, -0.152838261505772, 0.218719788507112, 
    0.449001266760464, -0.194542712859063, 0.105445103589155, 
    -0.0398613299644097, 0.244259287298288, -0.504545026259807, 
    0.0519319345849364, -0.422770041653452, -0.328223896063866, 
    0.0777556509466752, -0.390167024394012, 0.00988957277741517, 
    0.0426635284140858, 0.0547139036461406, 0.0545386892206841, 
    0.0553436136680868, 0.0548671896816517, 0.0422638062637121, 
    0.0214217534128923, 0.164377537086114, 0.154794080465295, 
    -0.0915644847910841, 0.0997309859393612, 0.600943655780906, 
    0.25934535296267, -0.213411242148624, 0.401436217284395, 
    0.537160547419877, 0.168708697200254, -0.0276334937022293, 
    -0.0296305260930374, 0.301847281393318, 0.402829115522303, 
    0.284326724661884, 0.228985646558343, 0.305916808972408, 
    0.345717373467662, 0.305587822151216, 0.251626395711555, 
    0.175506728832584, 0.320474632190058, 0.528551351878752, 
    0.281280722654701, 0.0624507047611875, -0.0410202240219414, 
    0.455011541550653, 0.276431083241534, 0.210505247590405, 
    0.542356471293659, 0.249204037787984, 0.101538459703871, 
    -0.464000930492121, 0.201563182658706, 0.534616460166219, 
    0.135208718384781, 0.827549024418699, 0.693241242993742, 
    -0.00141039711672253, -0.0444544415864328, 0.853472842927947, 
    0.477080934584481, 0.320927086678379, 0.710678137106176, 
    0.156948756247354, -0.0687068591858506, 0.493888802826428, 
    0.149035351402552, -0.244025177088503, 0.0907212136968812, 
    0.277862572359626, -0.132816811232527, -0.239416641902678, 
    0.129713885298511, -0.528910744271227, -0.125550128511995, 
    -0.208325616836719, -0.335179727553046, 0.0699864317889443, 
    -0.130779036645621, 0.080849989435922, -0.375397250776625, 
    -0.12035351624669, 0.130920298696283, 0.0985457452947919, 
    0.0359028691448895, 0.193750848327288, 0.171956596723977, 
    0.0431117888131602, 0.0359959534582377, 0.305249014535473, 
    0.129501516889146, 0.065441981821769, -0.00471809951822833, 
    0.523320586910315, 0.263447312208937, -0.0299149653891942, 
    0.65627931968575, 0.299203288216815, -0.0600265448921525, 
    0.122451426349342, 0.590823652097212, 0.228595414913876, 
    0.100410374180617, 0.0717160158900409, 0.0748627225614523, 
    0.0643687597159017, 0.0697168699507855, 0.0644984891566478, 
    0.0813911200896895, 0.0876525756142148, 0.0384615600483502, 
    0.0710102913995672, 0.11135207109406, 0.13444387577621, 
    0.141365761665766, 0.153065359041782, 0.151969354303539, 
    0.151597467330261, 0.174927842968884, 0.153080186793676, 
    0.113117411681977, 0.179727873581776, 0.215825070513557, 
    0.211573997165194, 0.223080395615478, 0.238789992680389, 
    0.216119031147104, 0.218281340696594, 0.286022713409198, 
    0.316719997608267, 0.30050106498035, 0.254584950341201, 
    0.171320132263026, 0.352230717755091, 0.502120099350686, 
    0.241843278315197, -0.0040466701218487, 0.507841954711342, 
    0.493515687029903, 0.126496910935959, 0.048688794012715, 
    0.761137762604917, 0.0872821516734156, -0.0775900497539443, 
    -0.171295485606984, 0.434079650753452, 0.395696730261722, 
    0.398013814606982, 0.441558305591337, 0.189177531258753, 
    -0.131351248880043, 0.690355578502421, 0.224891040448223, 
    -0.00349574747930269, -0.0148127613762233, -0.0538262713852215, 
    0.177883834643216, 0.0760538665165126, 0.724039400641328, 
    0.122455698857574, -0.129768116672085, -0.159384837986309, 
    -0.0720554994464634, -0.110940979593273, -0.0826233487011074, 
    -0.0162412280393904, -0.0515242394446456, -0.0299031085523585, 
    -0.0604307440995966, -0.114847559273538, -0.105810842708415, 
    0.00614492264530644, -0.00518619161146326, 0.029290810947345, 
    0.0122665654570966, 0.0408589311822694, -0.0150312409540503, 
    0.0297726017165102, 0.00837642994305786, 0.0485135359058596, 
    -0.12256685243854, 0.0572244497149407, 0.33704473806843, 
    0.226544628746728, 0.0804688401885415, 0.25507093991809, 
    0.166545622423763, 0.0245828883500601, 0.362700524458186, 
    0.364735080525827, 0.493464227915942, 0.444826719689307, 
    0.509102326602065, 0.870348123282101, -0.00382859570442134, 
    -0.103822089943137, -0.10640740847161, -0.0487442286212046, 
    1.36522754861499, -0.196035549348425, -0.0485035576099947, 
    -0.293984055531382, 0.0258603753005633, -0.2105231429316, 
    -0.125131306424955, -0.132008736643348, -0.139705582089873, 
    -0.0818091779258366, -0.169393641535005, -0.00411271671531421, 
    -0.141405239584055, 0.00833305941090064, 0.111522412140018, 
    0.188730973863846, 0.194816979253654, 0.140522457440149, 
    0.12935724800918, 0.221671346593524, 0.237082318109402, 
    0.206020606983367, 0.189341881498651, 0.16798889271608, 
    0.162210551705554, 0.161498302626777, 0.164130861341691, 
    0.171696509039748, 0.158961022659224, 0.147030828554518, 
    0.156545627841786, 0.170420872635605, 0.212550182420801, 
    0.200358935393566, 0.0506550364450328, 0.035183488117072, 
    0.400345366440091, 0.31753360040114, 0.141633775153999, 
    0.0848826854622747, 0.0715956554863967, 0.00481463660185805, 
    0.659349077544531, 0.448860418642945, -0.092098082800517, 
    0.622115903867964, 0.549898636024966, 0.0684504352986439, 
    0.295507815872952, 0.654552872876272, 0.367842603784804, 
    0.618484349085984, 0.601818102577305,
  -0.335018747363624, 0.583114607944967, 0.379267479583173, 
    -0.112095511736301, 0.214495500097885, 0.723090515690354, 
    0.139881759405673, 0.248973689458223, 0.977967595988622, 
    0.147471886596402, -0.0433725728940663, -0.00104850035637842, 
    -0.00815686732074956, -0.00700583793641538, -0.00759377052782324, 
    -0.00584104058281383, -0.00836448637015609, 0.0162367146149671, 
    0.112155356240414, -0.149206061311273, 0.286914045242707, 
    0.242837227707181, 0.117145428219995, -0.158332061622464, 
    0.309941141872133, 0.296332709682239, 0.0798451379531262, 
    0.442513766048232, 0.373796489164198, -0.107111767801366, 
    0.213190502700942, 0.538460028004998, 0.123092441967802, 
    0.114597652131042, 0.0655611748134638, 0.507100427901325, 
    0.0794039433273511, -0.124430726009449, 0.336598836084607, 
    0.193175718145754, -0.265331028215635, -0.0605172594016355, 
    -0.122608175106644, 0.0188346303189477, -0.135935328777487, 
    0.0320045604245957, -0.478249381142197, -0.0348087106362631, 
    -0.192680452628667, -0.206310629632596, -0.057902796761293, 
    0.0823393522875514, 0.145310210249809, 0.16419513751236, 
    0.14229791919982, 0.145669150728002, 0.204431105742112, 
    0.205375553996081, 0.135692213743844, 0.0983071978347368, 
    0.157203133684872, 0.190056517466154, 0.189127270886033, 
    0.221261474691682, 0.248007636740773, 0.203630521951705, 
    0.216560003009882, 0.285695804011637, 0.205039993832739, 
    0.228194386505103, 0.485789029679235, 0.246766713129067, 
    -0.171184133772839, 0.335772335707836, 0.504590918337173, 
    0.167654218551946, 0.0889787352448245, -0.216967713334876, 
    -0.117256754331008, 0.257644738045914, 0.607567922943254, 
    0.207492972021103, -0.143964063613086, 0.134840456221895, 
    0.617487837869732, -0.0248898401954751, 0.245901757233312, 
    0.728530819886608, 0.199680249681428, 0.0509115898865254, 
    -0.0572492019956321, -0.16985979929549, 0.224300443415526, 
    -0.0798410990065955, 0.171674261321427, -0.186345259438044, 
    0.108641039792214, -0.184914899697279, 0.0618029162030785, 
    -0.227626951067367, -0.0203821750494762, 0.0740800344279556, 
    0.141314229680699, 0.186792168463325, 0.201448169912381, 
    0.18604261357017, 0.223454720475049, 0.279000728573272, 
    0.239380709136434, 0.219052098020659, 0.279581560460986, 
    0.201999785936121, 0.135365673929928, 0.391664867398629, 
    0.42443410407537, 0.185012024813793, 0.0432311640655314, 
    0.26433455999412, 0.429101689902218, 0.49584450542812, 0.295174106042062, 
    -0.0249829953227626, 0.124452350120234, 0.784537222779363, 
    0.0535935497369273, 0.00418491638840682, -0.0533927246016158, 
    -0.0790987929401408, 0.0824071018336125, 0.815751977109835, 
    0.313521784140599, 0.0727389586299867, 0.389985751901904, 
    0.0104163413378835, -0.233418852572069, -0.347196183207097, 
    -0.160230257368976, 0.513918745064857, -0.0759468690877352, 
    0.101580654470716, -0.376589401025773, -0.164411771541855, 
    -0.168131196437307, -0.281020866848139, -0.14210701950434, 
    -0.234298015440496, -0.202592324313909, -0.160674512523442, 
    -0.138208822116924, -0.200853468980788, 0.00355711648453359, 
    0.0824526570393221, 0.0302965560026345, 0.0284521694912254, 
    0.0821135403567848, 0.0756248809731818, 0.0993340808894532, 
    0.0622735023466984, 0.0454882654637487, 0.0998390932399748, 
    0.213139703548331, 0.0653794793433738, 0.0337216689937595, 
    0.449645910221586, 0.228022413433198, 0.102650312189714, 
    -0.0459920135735281, 0.253527397746641, 0.247248911498439, 
    0.328144113168713, 0.415614174455372, -0.340874383948365, 
    0.486741885588904, 0.90118099814305, 0.0188061644163101, 
    -0.0536854521078416, -0.0975214596291543, 0.43994207161019, 
    0.833269476321483, 0.0332070756501123, -0.0568284904674398, 
    -0.0798473716636667, 0.0747908633529751, -0.0327131189285388, 
    0.0530357019668198, -0.0669277588064078, 0.0226899771991662, 
    -0.0131479667556893, 0.0489284493065438, -0.0857487758346247, 
    0.038041304334178, 0.104044478287272, 0.204472050232375, 
    0.188116904195764, 0.119898878378347, 0.235264325686357, 
    0.397148326436354, 0.30966357961992, 0.171153079664203, 0.13388971542666, 
    0.297027364704438, 0.387485015143415, 0.331473048736932, 
    0.311755311210189, 0.315472038526323, 0.242526001932916, 
    0.214399612384294, 0.339878856596146, 0.319215019574761, 
    0.162237410252781, 0.105759116682193, 0.381760786618839, 
    0.422701622248585, 0.142103474121015, -0.103752369242683, 
    0.0978935625420446, 0.567057612847096, 0.071294863517291, 
    0.0603608082680239, -0.218428421141882, 0.368486997093861, 
    0.321627252798382, 0.132337510916098, 0.118137803833545, 
    -0.166500513751411, 0.596557021109544, 0.0972719108495581, 
    -0.205956851023313, 0.406403867488629, 0.127870292295175, 
    -0.283564870436819, -0.0511210069448662, -0.0801587952893351, 
    -0.0164897751530036, -0.122731245701383, -0.00231994279882218, 
    -0.124084336898554, -0.146081558420545, -0.153106015789618, 
    -0.0913611077450272, -0.142654297405466, -0.222995966524433, 
    0.0859720808578777, -0.0628327855752878, 0.0755394631438069, 
    -0.106148952680972, 0.00114624732152231, -0.153610580894779, 
    -0.0257399209385632, -0.218344328938993, -0.104415601571333, 
    0.0555707635561325, 0.0968078348895925, 0.0412025588747487, 
    0.0152028138134044, 0.0671474029290218, 0.137611816389028, 
    0.272616636088071, 0.220261803793522, 0.0928858900136894, 
    0.727868044389587, 0.0990261381850381, 0.0459242415014945, 
    -0.329481839735386, 0.0715337310877277, 0.720859193218485, 
    0.129584774770574, -0.159969450372946, -0.020187130976998, 
    0.535687640149945, 0.196799489693075, 0.107822456053926, 
    0.128055211296687, -0.266916553021319, 0.368404726660686, 
    0.393109371805556, 0.140844282647863, -0.233958713213143, 
    0.209887181648942, 0.394275672115578, 0.0326467421326288, 
    0.00316419120390995, -0.0957135120193843, -0.0880865429547789, 
    -0.0887275146134585, -0.0576605850837914, -0.0116894012441594, 
    0.0207314456606952, -0.112504239804982, -0.140075619312932, 
    0.054759251302742, -0.070278358188518, 0.057218015335688, 
    -0.05469875174193, 0.0425088024901078, -0.0969974214396643, 
    0.017133855708449, -0.0705982153631695, -0.029187505177643, 
    0.0508766433045365, -0.101375390379834, 0.199315835059493, 
    0.149542411200015, -0.0326265897127842, 0.0441459212953641, 
    0.343648887794333, 0.0554237463135273, -0.0354673350516739, 
    -0.143929286077239, 0.00522627047355132, 0.648984599344804, 
    0.163800303619502, 0.0450912698082496, -0.554787696454769, 
    0.200215815810165, 0.554787251852909, 0.620667500667913, 
    0.438500432662589, -0.286652102801669, -0.619316301855887, 
    -0.402804398290431, -0.291612476363806, -0.00618384793489508, 
    -0.419296042456301, -0.0802802176799536, -0.22290844478801, 
    -0.217979892688298, -0.0134974588530366, -0.406975102733993, 
    -0.0231669194643818, -0.108440749495492, 0.016851040436723, 
    -0.238230407937195, -0.0490604277815937, -0.326262964799718, 
    -0.194726230153033, -0.0563775995127881, 0.150418456457849, 
    0.0300519112222154, -0.265328202761915, -0.00599023846522408, 
    -0.225105148164955, -0.186457657043121, -0.0685670366076505, 
    -0.209194410874352, -0.0659554421192986, -0.210259307081588, 
    -0.118517411006822, -0.0462024157857709, -0.116939876344088, 
    0.470294986838894, 0.0478179204669503, 0.116280776480415, 
    0.553771256648822, 0.0709469258533489, -0.0275222314534181, 
    0.0803512997936462, 0.387647756069334, 0.113746259030212, 
    0.154740144790497,
  0.174679704387622, 0.123512439659317, 0.16820395301068, 0.13522536544888, 
    0.151415271591156, 0.115475192159378, 0.0924743190844728, 
    0.243563033486325, 0.183718365372135, -0.0128175338530853, 
    -0.0589027126119809, 0.0755842278362153, 0.598732746763873, 
    0.170672640211433, -0.0962410150095621, -0.0843117113407884, 
    0.470495357207509, 0.294336663556829, 0.0989105018894242, 
    -0.0937333468609082, 0.0301880231465137, 0.496471739462827, 
    0.152567028584459, -0.0966762987763005, 0.239848499778758, 
    0.272438798815268, 0.0454160612778634, 0.41748793364389, 
    0.293668067848089, -0.0210341575947145, -0.0967409100695476, 
    -0.0359728973135921, -0.0595658536174151, -0.0690672312458525, 
    -0.0122540494434225, -0.075890266237094, -0.0308621357475641, 
    -0.00659334808277409, 0.0289412196399313, -0.0970481953075817, 
    -0.0238371347530534, 0.102496924323878, 0.152881913032689, 
    0.254226276223867, 0.204479318516759, 0.0723037129278546, 
    0.362146226748719, 0.192059573247757, -0.197127545334033, 
    -0.100242557574374, -0.350817297743735, 0.373762904417998, 
    0.0863255467466599, 0.589253247325115, 0.962112110687466, 
    0.284551867236346, 0.118140766657859, -0.147683455066999, 
    0.229237830404284, 0.594805280376766, -0.129040376072877, 
    -0.000573663056678622, -0.213576314773415, -0.07542466987496, 
    -0.0169740357611176, -0.151857719499294, -0.0310573659221798, 
    0.0122381416961984, 0.0384115115053704, -0.138931435020466, 
    0.00825174967084098, 0.0883979614947257, 0.190232085745023, 
    0.217490751002723, 0.2354661626507, 0.29000707112973, 0.25351115602281, 
    0.155046698796719, 0.175600990259464, 0.339707906870787, 
    0.349419064836536, 0.268143393873623, 0.216291052322078, 
    0.20766396894484, 0.209862330269753, 0.189888687085553, 
    0.181063675236274, 0.186525691987264, 0.169223253857072, 
    0.211672609923761, 0.310828377114036, 0.182621736848351, 
    -0.0588082942756411, 0.347219825825745, 0.386859948475237, 
    0.0993105381741601, -0.0220533893650727, -0.103779435852152, 
    0.586400028343495, 0.21576285948723, -0.164752905223329, 
    0.260119963240312, 0.469762013131725, 0.118951702734266, 
    0.0330444229947779, 0.530453613263946, 0.0726050872201673, 
    -0.428363806177593, 0.0751842823913949, 0.444721167741778, 
    -0.323590240996336, -0.0954593519935183, -0.163435578421088, 
    -0.0970847274450235, -0.158338651381872, -0.12237108704021, 
    -0.101624614368764, -0.111859814554209, -0.15363702993381, 
    -0.0595523079377948, -0.00152263653162532, 0.110150600893351, 
    0.0328293937522721, 0.0866132888198156, 0.0223056349647042, 
    0.0722209833175584, -0.0476746845758442, 0.0290336729287515, 
    -0.0130660274034985, -0.0245577651463052, 0.0332371640963225, 
    0.0648552501331507, 0.0801807931375558, 0.097877761909376, 
    0.107480521952392, 0.0743460367958073, 0.101780277337399, 
    0.183074758954374, 0.0453366073526803, -0.13480559548686, 
    0.148050930397585, 0.380121629124472, 0.0447797690118777, 
    0.0343325198191093, -0.28737430587937, 0.793050120568768, 
    0.191883101114189, -0.18829831872606, -0.112890751310205, 
    0.55110833118337, 0.67409323281007, 0.296822183371994, 
    0.0121567684570039, 0.465786911802068, 0.337779185561271, 
    0.0799500101210213, -0.430212714463706, 0.352499983900932, 
    0.393519007334127, -0.093594225042644, -0.117884938255868, 
    -0.227233206920624, 0.0657321145209815, -0.128835936476707, 
    -0.0123644999476734, -0.0937336669750283, 0.00837329269822124, 
    -0.124742108759076, -0.0414370494016936, -0.0782080563447757, 
    -0.225590773337506, 0.215713946781254, 0.325696390864591, 
    0.0862377860686316, -0.149340844221103, 0.565551143452849, 
    0.321318708462449, 0.0613823791814962, -0.0298856456320551, 
    -0.17869830012918, 0.0963422278043224, 0.420562445132493, 
    0.384998943145165, 0.377270454238565, 0.48237855161626, 
    0.390385812863529, 0.195715036333217, 0.152776171261263, 
    0.461900647105927, 0.41465440936591, 0.163434046060707, 
    0.174016066864399, 0.408858410974819, 0.277083822391488, 
    0.100385122770791, -0.116454627145673, 0.303890245279788, 
    0.339362429902635, 0.158095758670089, 0.141996135049018, 
    -0.299856562895027, 0.191199516999496, 0.355378197288972, 
    0.0760482718963819, 0.675196243034286, 0.482009421597744, 
    0.100303535844897, 0.148984517395142, -0.350397571492813, 
    0.207440882722669, 0.426854803761872, 0.0555781296403942, 
    -0.212527385788719, 0.00720392986274231, 0.413050386904421, 
    0.205470341937906, 0.0689751725338645, -0.156716563998844, 
    0.27532073072796, 0.164398136355127, -0.312287276763961, 
    -0.207381115864369, -0.117753976927299, -0.234161280769023, 
    -0.0966565188658284, -0.223070033410551, -0.117353254426749, 
    -0.198180741379533, -0.00387974873849348, -0.257069736202354, 
    0.0164946478677954, -0.0201133042046865, 0.0303332989919175, 
    -0.0889255366966122, 0.0372070548427983, -0.11232331438712, 
    -0.0235572848965864, -0.0226044601620217, 0.0506348746418917, 
    -0.0957623099909671, 0.0559932306883041, -0.00134657177427862, 
    0.00357832865225012, 0.0201108582790192, 0.0256033714643336, 
    0.00937365201427598, -0.0110828103677571, 0.0502810135051565, 
    0.0221853289338983, -0.0199364823113195, -0.0739964131080377, 
    0.029454744050086, 0.378403346350404, 0.159612897517178, 
    -0.0109980440349214, -0.0273344279564394, 0.0997057978344635, 
    0.516075711237582, 0.357211062381358, -0.111451047796787, 
    0.640789635722233, 0.375957700999053, -0.0239356636535322, 
    -0.118152032429821, -0.272399059098055, 0.515294399376912, 
    0.225019713280875, 0.489230778275069, 0.97758573111334, 
    0.181061609530517, -0.106897061489998, -0.146893999196637, 
    -0.0712422224747821, 0.150526730422682, 0.139440864746451, 
    0.114735272997301, 0.0844069989625273, -0.0477412526866335, 
    0.194989684758326, -0.0996438292746516, -0.33148290093657, 
    0.086341843510996, -0.22952951422859, 0.0262486389559552, 
    -0.224459886909793, -0.0306200860134764, -0.153791264582081, 
    -0.00585251401024782, -0.226168171364902, -0.0422258348294373, 
    -0.0335274737383841, 0.0738363367525369, 0.0397578002580962, 
    0.0700581379796724, 0.0295612345990483, 0.0757495239139026, 
    -0.0262922890244588, 0.042414179387568, -0.0416643134368223, 
    -0.0201160905285945, 0.0393719969912596, 0.0551103854071839, 
    0.0827136661913186, 0.0597749607903193, 0.065562638373762, 
    0.0616662912550379, 0.0662547845546118, 0.0912332906171864, 
    0.0789758815385328, 0.0234097967589346, 0.0696440555213457, 
    0.131064932195805, 0.210489772801784, 0.180063421109747, 
    0.0714708019253824, 0.154358162258838, 0.380555263484774, 
    0.191951737443815, 0.0709595745969952, -0.0650093157351677, 
    0.571129685859148, 0.152890633162017, 0.0443191516853606, 
    -0.2491869035322, 0.0594375573317183, 0.633724037083426, 
    0.0927519345015367, -0.224422694870254, 0.158397456923969, 
    0.525717261247691, -0.0557811506571641, 0.0186257132711902, 
    -0.199118830695855, -0.0675845362108858, 0.077895412697263, 
    0.3599218233795, 0.210492743729555, -0.113624710389781, 
    -0.246680162256557, 0.0530880528282912, -0.212397031708901, 
    -0.0757706241060468, 0.160264252057302, -0.501164124052073, 
    -0.0170636636312918, -0.12623298168579, -0.0327344808809276, 
    -0.0095877486550932, 0.0924879000829177, -0.289878679894856, 
    -0.0133303700823163, 0.190474653854265, 0.130061594059099, 
    0.125737495961359, 0.293402768289584, 0.237523551442148, 
    0.0899582794806248, 0.129466688023543, 0.374831518034615, 
    0.318209851319761,
  -0.0549480696208561, -0.0959820356344107, 0.0595264582762465, 
    -0.0975414010174066, 0.0139822012526089, -0.125013333033514, 
    -0.0179972780758113, -0.108830314722508, -0.0570046740310734, 
    -0.0407556879202733, -0.0130285703110239, -0.0220776898453172, 
    0.203116862872385, 0.325821027956514, 0.182380536305645, 
    -0.156420300997787, 0.174740475087496, 0.373650240029491, 
    0.33208272670139, 0.254234303719673, -0.423794416732858, 
    0.680372888143348, 0.89544199092345, 0.225998323654339, 
    -0.327755030394696, 0.278930763598762, 0.719264003725541, 
    0.315120322499537, 0.126771787544915, 0.194453016587594, 0.4805810165038, 
    -0.205763290048962, -0.202233783332028, -0.0551470217745251, 
    0.216984396072733, 0.20117985713717, 0.131929460181424, 
    -0.151080225702864, 0.178194569461495, 0.0777754142986973, 
    -0.107178227395829, -0.0635463321006479, -0.139536161838573, 
    -0.125178500477254, -0.0865195388828441, -0.078432191619923, 
    -0.109711743989653, 0.0305405193968043, -0.165413790745515, 
    -0.0343661798532485, -0.137540835928844, -0.0848012375897205, 
    -0.0628931802989448, -0.115140986492957, -0.0313956291633614, 
    -0.11019194674171, -0.0120185629192661, -0.0971730650515426, 
    0.0167604783654031, -0.100740915346785, 0.00884880828722694, 
    0.0440018436866943, 0.0523103462550136, 0.0516953402955339, 
    0.0523081282638766, 0.0588044787182722, 0.0690939252554847, 
    0.0612191369137466, -0.111031551013753, 0.112298958263068, 
    0.488195166868831, -0.0109010926922279, 0.19812872993351, 
    0.6064057078187, 0.115162846925992, -0.0538328148796185, 
    0.260115350775639, 0.374200209494277, 0.0172560623948923, 
    -0.259372452311739, 0.349119706943765, 0.471491939205809, 
    0.164702101120052, 0.0410284042379149, 0.242345726630963, 
    0.197087561012923, -0.0478210247622515, 0.279136108616098, 
    0.314705695052695, -0.0588488215403831, -0.119510323531793, 
    -0.130492488659189, 0.0162697989649444, -0.121071071759004, 
    0.0316732061776146, -0.189738579594235, -0.00290229727784756, 
    -0.201010270431034, -0.11367497955684, -0.00882718784018464, 
    -0.0947989600570616, 0.0822748640376221, 0.205716879385759, 
    0.0563340329342855, -0.018332141759586, 0.077636613240536, 
    0.186429086684698, 0.15922594283253, 0.226331210188498, 
    0.569262891614465, 0.0848862698462508, -0.21530640870184, 
    -0.111861344709777, 0.690651650157848, -0.121529539229046, 
    -0.0234309688534007, -0.126381048161257, 0.961947467776995, 
    0.0651330698030102, 0.0388102441972779, -0.213296398561559, 
    -0.159015997940688, -0.131822442034378, -0.0858504169896823, 
    -0.213384174124976, -0.108860590869464, -0.0104482062804905, 
    -0.249161259380621, 0.111038814362192, -0.141972363420139, 
    0.0624608748914496, 0.0554043722007024, 0.121194669740413, 
    -0.0788980399725412, 0.0279328127606354, 0.0376653142819481, 
    0.086349216826504, -0.102437389192782, 0.0652595020559991, 
    -0.0219586739234149, 0.0575807591184926, -0.0542128261105003, 
    0.0108816717211417, -0.0332348867392919, -0.00533990527851594, 
    -0.0584050911628729, -0.0351191603038074, 0.0101177618417332, 
    0.0519248913313155, -0.0784572078917475, 0.0664039945085464, 
    0.111746522137767, 0.0682289403300606, 0.0699699788043287, 
    0.0600262980380326, 0.154879143598258, 0.226188282108079, 
    0.0733759015614977, -0.00530320440763907, 0.0473406096327441, 
    0.110673727448081, -0.238185325434758, 0.523538912215004, 
    0.29325957384361, -0.134219892845057, -0.0581003478102106, 
    0.788670364335064, 0.471053865088338, 0.241469743971287, 
    0.344209057388324, 0.120154788708288, 0.381730463902348, 
    0.712674401523928, 0.156955075900658, -0.177943589829868, 
    0.24645641849068, 0.237148492183881, 0.277716114926643, 
    0.687791577949463, 0.281456201214598, -0.0347250898772344, 
    -0.00727917166966739, -0.146340800925084, -0.0305854504767763, 
    -0.0626866159077487, -0.110729270644828, -0.0414331652941052, 
    -0.16309486155329, -0.0547244810178057, -0.0495816840521132, 
    0.0224274024299737, 0.034931416519601, 0.00708796840417561, 
    -0.0063522767650273, 0.00591994975168925, -0.0199103385341176, 
    0.0312317024606719, -0.0276255500485676, 0.0201485805006602, 
    0.0609229822946236, 0.0301356223102845, 0.0692478843181945, 
    -0.127003897921351, 0.062866415514884, -0.077255869985246, 
    0.0259733796158073, -0.173037672675532, -0.0333777516361033, 
    -0.104198567988491, -0.146401603265326, 0.0184362558986864, 
    0.0641065504614928, 0.0218559491359084, 0.0709964997571419, 
    0.143855011747971, 0.0889342386780977, 0.063414060747702, 
    0.0747691176589112, -0.0770791497649482, -0.0322102070137166, 
    0.435580005753187, 0.303159261194438, 0.247412178906706, 
    -0.29892166627423, 0.54249224907515, 0.478252408318368, 
    0.0722292495678626, -0.263402277604047, 0.0976378595556786, 
    0.568282257908949, 0.024055845602709, 0.0051938745773222, 
    0.133896870869373, -0.226399448985917, 0.395160478353641, 
    0.297231546723247, 0.324709702046294, 0.207938670766901, 
    -0.248749292486652, -0.142447606363233, -0.193557829223296, 
    -0.235159443418161, -0.146088966605703, -0.287045103237263, 
    -0.0946767160421898, -0.298259953741906, -0.125039492282464, 
    -0.228936404113734, -0.108608813384673, -0.193725408446959, 
    -0.0177793211603251, 0.0261006631902669, 0.0139310707781466, 
    -0.0213593936168975, 0.0956628347126883, 0.0297698254739422, 
    0.069265235284175, 0.0400014415693598, 0.0579683393980238, 
    -0.0230401725936358, 0.0524917322061811, 0.0462832927355289, 
    0.090204933625175, 0.202855906368078, 0.116320190668065, 
    -0.0141960173395988, 0.18387749536048, 0.174706640982876, 
    -0.0297107991101833, -0.00453907799413679, 0.294878233088779, 
    0.0952268252183212, -0.241449859615163, 0.184079189638922, 
    0.418811680862452, 0.183601298346833, -0.273160030655032, 
    0.397057623613662, 1.27284608567477, -0.0430742418606121, 
    -0.33258097764011, -0.177380576014945, -0.079911171142513, 
    -0.186360735190405, -0.104915176163657, -0.0953173260334964, 
    -0.307903504526261, -0.16923298695311, -0.380374134081721, 
    -0.340911542333183, -0.194911686119353, -0.163920814523868, 
    -0.0246610137195459, -0.0665730098231154, 0.368713820231261, 
    -0.207270104322618, 0.0911821409218117, -0.076527115408888, 
    0.0567389251994583, -0.4332393762299, 0.0268087250580551, 
    -0.0960238906550144, -0.0706715061781606, -0.0548608886340915, 
    -0.00039154828545436, -0.0238988430046892, 0.0100147007542866, 
    -0.00404185615078775, 0.0313372728612144, -0.213879519291976, 
    0.545322944001365, 0.174264385382945, 0.504787932425451, 
    0.434168384813908, -0.306443276707174, 0.19384247291409, 
    0.893857690457268, -0.0651262333781754, -0.193719552800096, 
    -0.111572375159084, 0.59659916921531, 0.352339291798402, 
    0.128135117744458, 0.0159340322965756, 0.196449648658807, 
    0.335813475019929, 0.348339432778821, 0.248618563913516, 
    0.0485022056948866, 0.267764065852278, 0.583986868024878, 
    0.320955712107965, 0.118277751735942, 0.228264389455487, 
    0.313758260829445, 0.129790747581646, 0.00689820753164919, 
    0.23092397044603, 0.366720827444403, 0.0855743681103015, 
    0.00582827591392709, -0.226321089812564, 0.169123434107715, 
    0.593633349123979, 0.15555046154441, -0.175808530868352, 
    0.0960208863315132, 0.398389796423643, 0.160752046349501, 
    0.176514578645107, 0.426716202977423, 0.224792220485432, 
    0.0267036887578364, 0.264090175976457, 0.364483164010617, 
    0.0452289630925845, -0.200914383642803, 0.145264723866964, 
    0.201029092516913, 0.0138732990146516,
  0.39276572534717, 0.300754754635674, 0.197289411657177, -0.320669038375977, 
    0.177806192655538, 0.503564111536835, 0.0181175059435747, 
    -0.101405471040903, 0.22948553555246, 0.515107324727346, 
    -0.268364391233543, -0.144760233813584, 0.1117316078858, 
    -0.125811604138882, -0.0277413095010303, -0.175086769760382, 
    -0.0152467206924514, -0.024018717684862, -0.0941054937110834, 
    -0.0507494373600908, 0.00448874656602197, -0.12000660457206, 
    0.0734459352046929, -0.0503278485812904, 0.0795075749318841, 
    -0.131156351931525, 0.127036682175612, -0.260534976090099, 
    0.023872861916898, -0.169525695498603, 0.0195322616728231, 
    -0.0420194625085074, 0.131983747083413, 0.200879665947042, 
    0.070470257929375, -0.0315464521209216, -0.0551751006138931, 
    0.36266372474467, 0.106443601786879, -0.0263947596523099, 
    -0.106170016672011, 0.67063290322991, 0.50019136210436, 
    0.322268388949664, -0.20619490486447, 0.495434476966284, 
    0.518930506484211, 0.197729997389079, 0.0825964676055394, 
    0.807394260051261, 0.405531842019269, 0.159439765560089, 
    0.033102337458137, 0.170524616561038, -0.221036408570835, 
    0.593942374151903, 0.494721286407282, 0.185207594982786, 
    0.752434996460012, 0.460724477670956, -0.0816115037821154, 
    -0.23912285872185, 0.206855668037855, 0.107484968669976, 
    -0.174346400346256, -0.016965770201343, -0.103670865118652, 
    0.148610952967195, 0.0363503766077535, -0.18889936130561, 
    -0.135551084053271, 0.0521510928948165, -0.17770623395025, 
    -0.0204068223978744, -0.140209639206274, -0.0904394954872822, 
    -0.0712716250474593, -0.0783950158109676, -0.0773592898599595, 
    -0.0301190303816859, 0.135673964415637, 0.0356926246937678, 
    0.414021608848536, 0.167233907203894, 0.0590243989478045, 
    -0.108074636499002, 0.231283434831774, 0.225747251126741, 
    0.202189251622567, 0.418299702905084, 0.336478631772363, 
    0.0379176032522592, -0.312525782329158, -0.192993498424878, 
    0.627267626809704, 0.390899961268946, 0.156102628898623, 
    0.43113339790518, 0.364603213842071, -0.0499263822396791, 
    0.329128723272968, 0.65509921166656, 0.337400603228778, 
    0.127647942882112, -0.125511534568816, 0.224278121556359, 
    0.224641762321391, 0.0675411957852772, -0.110018115994021, 
    0.133453164734869, 0.199921270383934, 0.0483802091398558, 
    -0.00552299076315656, 0.00127941385677632, 0.0632925413521243, 
    -0.151532938242581, 0.0226446091294806, 0.121203378555671, 
    0.0311034027637234, 0.0165006378717467, 0.132523461381516, 
    0.0410242879597135, 0.0214689306741037, 0.0205091350835879, 
    0.0156604834512052, 0.0265384137888407, 0.0859163634206637, 
    0.0314534289005091, 0.0236132620915858, 0.013363001818004, 
    -0.00891752785682948, -0.0770803548172761, 0.00865252471549352, 
    -0.0128455503003727, 0.0184114158376783, 0.014850586919618, 
    0.0695700025861132, 0.0202044927182128, 0.121340472566701, 
    -0.0844413605796085, 0.14340408956107, 0.244302141845877, 
    0.123875355363371, -0.054931367637334, 0.17218214101597, 
    0.0675763297978366, 0.443293747849735, 0.434815104680004, 
    -0.069234329725246, 0.0120539110839691, -0.120987105386406, 
    0.671960745746208, 0.54056549213592, 0.451631804552198, 
    -0.361298134767995, 0.487760407487258, 0.478603905081963, 
    0.125434980798058, 0.123923231775036, 0.165447876383492, 
    0.594998048964421, 0.661903280022626, 0.141251702626769, 
    -0.0225634443937285, -0.0161050971696526, 0.249618400305493, 
    -0.321492126097636, 0.399712100008646, 0.262687090026796, 
    -0.190200213459407, -0.0972728445475529, -0.165452627090689, 
    0.148673972620174, -0.213669818383457, 0.00131447920966246, 
    -0.128609444850865, -0.0783931166463307, -0.131630344181548, 
    -0.215734160012272, -0.0650648351440021, -0.101597707639091, 
    -0.0750113677624171, 0.0836520338566168, -0.129802252631065, 
    0.0579378231067972, -0.0417386810473442, 0.00945693758435465, 
    -0.0157845342810848, 0.0519493085550723, -0.139690596655099, 
    0.0793745542858873, 0.112866368457727, -0.015087853864687, 
    0.111184076356245, 0.352701941678114, 0.187232704329998, 
    0.0251526413096932, -0.0590463592972958, -0.212868466784991, 
    0.251209588099651, 0.543769081699527, 0.234532021869804, 
    -0.275673966875199, 0.264594972744933, 0.550764484520079, 
    0.154596355535995, 0.0209993761633787, 0.221768835232209, 
    -0.268454452727453, 0.280546425329882, 0.789340460743667, 
    -0.0705948471166351, -0.0987990000655038, -0.246565816517783, 
    0.501079990104559, 0.429550819485283, 0.240121234721152, 
    -0.219862426189149, 0.357878731466055, 0.358738298610585, 
    0.0479587878563978, -0.011927214808186, 0.336184701639607, 
    0.553250053926351, 0.199062611098491, -0.133124753574117, 
    0.146415899813078, 0.411155740619006, 0.225039893619158, 
    0.129723108907162, 0.147114470947525, 0.071535542820603, 
    -0.11446724303129, 0.290321816516176, 0.455488472639691, 
    0.133582764856064, -0.0142619307099016, 0.177394555819119, 
    0.15605485729084, -0.0370311111348478, -0.0777576221128271, 
    -0.0600355065124169, -0.0774077932767137, -0.0741492474516542, 
    -0.0340934569718679, -0.0814155206077302, -0.00140267285614329, 
    -0.0641416709131932, 0.0433179164388411, -0.0953152415128367, 
    0.0768712262263602, 0.0330631638918997, 0.122128316692585, 
    0.363153667299686, 0.160299604383853, -0.1198871485121, 
    0.162820093761855, 0.380305114478287, 0.160432862353786, 
    0.0893086370616799, -0.16892035246184, -0.191036435028167, 
    0.388442205793112, 0.49615536738082, 0.166727749918294, 
    -0.195735099583584, 0.0246934181587839, 0.457465374695638, 
    0.314666939956894, 0.238315920681659, 0.337551951801036, 
    0.218813770692809, 0.0783160662639522, 0.0213794515019045, 
    0.00777808672135623, 0.174829757603288, 0.252043598407657, 
    -0.238842793174003, -0.141397309561204, -0.167887268381933, 
    0.0793525627988606, -0.174570939603472, 0.137521199391748, 
    -0.11993643007911, 0.150332202938787, -0.186523583508255, 
    0.109882456183571, -0.128332698862297, 0.122309858954609, 
    -0.196880884238603, 0.0871415136165545, 0.0242493565727726, 
    0.04507316082433, 0.0459111867622677, 0.0636625879799942, 
    0.035290559863107, 0.0682964900808646, 0.0473865786229419, 
    0.0580256031930722, -0.0206231831389364, 0.0415255878642839, 
    0.120317981920543, 0.0799358075621171, 0.0635400666429405, 
    0.244328161872852, 0.157766009666863, -0.0224278983140781, 
    0.306102105175858, 0.169772400405847, -0.0747653142463659, 
    0.106530697301768, 0.272249547392181, -0.0193200335349787, 
    0.859220383873327, 0.386772217778356, 0.0145629887290452, 
    -0.00308183945406057, 0.123556811080263, 0.185492286022183, 
    -0.172375587519218, 0.507249489041564, 0.381136117885465, 
    0.0109664551219928, -0.0330226633656831, -0.0365233100672464, 
    -0.0889887432087038, 0.121475995096912, 0.0701208404520724, 
    0.0905342541449644, 0.0795652925037787, -0.0942271717354249, 
    -0.0497316484476102, -0.308483466368729, -0.0667448897487599, 
    -0.192838521472432, -0.27904364121945, 0.0186253306270729, 
    -0.0451294704473412, 0.0699361336944818, -0.208238263235297, 
    0.0216088857682764, 0.056683143877611, 0.0578632065319393, 
    0.0796318783220071, 0.0845420455135803, 0.0570253377218532, 
    0.0639760724355226, 0.0987451412329868, 0.0750192480591259, 
    -0.00576902521415026, 0.135839604384763, 0.185904598496485, 
    0.0870299829386359, 0.0955662877147732, 0.301228309276485, 
    0.312941187765994, 0.185727232285605, 0.0867809229114299, 
    -0.122440972443109, 0.33348631114628,
  -0.281935415326587, 0.0192687459860778, -0.284027025118228, 
    -0.142809637754338, -0.107696957967648, -0.190037184606119, 
    0.00167356812146252, -0.128472037430432, 0.0885234451742136, 
    -0.230372747748414, -0.00222667589908017, 0.0849886607784261, 
    0.135475966722493, 0.168593785151047, 0.16930734794408, 
    0.113947037895632, 0.0922552816988678, 0.247481009137452, 
    0.193258289673271, -0.124536684605934, 0.294624832622015, 
    0.383669872662189, 0.0687190990722134, 0.361589408019889, 
    0.559968433228019, -0.0445015294601207, -0.195340452263534, 
    0.0617439428207586, 0.542089038961205, 0.0101838894924456, 
    -0.447535535419792, 0.0375291986989329, 0.595727945004655, 
    0.907627501673235, 0.213076387575312, -0.315539343974542, 
    0.121885905400512, -0.647084831814083, 0.426455281037979, 
    0.385302740767151, 0.049386816684268, 0.0765628952489363, 
    -0.169582966138168, -0.127110687896913, -0.0809541504144263, 
    -0.148643970505308, -0.0442698041810796, -0.158011057464744, 
    -0.091616607578093, -0.062277808045247, 0.0697911391376188, 
    0.0751291924888914, 0.0880217342696835, 0.089166398654208, 
    0.0508404541034811, 0.0997937555771069, 0.107852440635563, 
    0.101423672880016, 0.0813432258256255, -0.0305680482224662, 
    0.0800763684617993, 0.255404175775308, 0.195300879049805, 
    0.0866114773606274, 0.00075520255926137, 0.258455809402929, 
    0.294457549411814, 0.138635314793224, 0.0728746299067603, 
    0.227153953006793, 0.237953058017583, 0.167145351842403, 
    0.12117636571514, 0.117604837720774, 0.137740870856054, 
    0.124785529965025, 0.105357254915795, 0.133347195910795, 
    0.102783950907755, 0.03927355386484, 0.0816664269759719, 
    0.225758309528337, 0.203864276598567, 0.0664182478103816, 
    0.103620775998839, 0.398688883809929, 0.307973728002547, 
    0.0977961279627045, -0.212491150926064, 0.134867370461131, 
    0.540887931551177, 0.140273190134571, -0.00093923589580644, 
    0.0751000123977101, -0.174734266789881, 0.360585553737625, 
    0.687269571878732, 0.217715739057826, -0.284678552431416, 
    0.513618674898921, 0.492218362494882, -0.00989458852677201, 
    -0.100665740267334, -0.173979829977197, 0.221359236627078, 
    0.356460026149848, 0.0638385643709031, 0.448751789270939, 
    0.566048352831896, -0.124786634455182, -0.143776867312982, 
    -0.113400330086404, -0.0517335897408632, -0.114937790128358, 
    -0.147554105072224, -0.104865325231249, -0.0302617973213096, 
    -0.197939951213895, -0.10136333035601, -0.19387136254415, 
    -0.0161484996209478, -0.184273828297774, 0.0675827254524069, 
    -0.0401944556109298, 0.0698108011174883, -0.151087734201434, 
    0.0255137320048644, -0.112236507094117, 0.0264693390380711, 
    -0.200386385863695, -0.0124354728164252, 0.0426953058597551, 
    0.0640197866558149, 0.108982476992598, 0.143589274417035, 
    0.113696619696771, 0.106849967264936, 0.170853811559139, 
    0.11806139335996, -0.0347764155770837, 0.192491048801474, 
    0.338619927269086, 0.140606360339821, 0.00988093674582892, 
    0.491672850763241, 0.359281303599914, 0.100701973992022, 
    -0.154625749980856, 0.215160218269188, 0.438886044982475, 
    0.365340283572226, 0.215904903470564, -0.203314783536584, 
    0.404279934161923, 0.404645846886902, 0.131238869567135, 
    0.0368334813781219, -0.173491421488038, -0.00120860208597756, 
    0.497265610160254, 0.349897480464347, 0.197905311802204, 
    0.0884910346288498, 0.00105302290210159, 0.0076928009100726, 
    -0.00669681098903278, 0.590422684367405, -0.0493691333849517, 
    -0.0344280147785171, 0.0280845354978681, -0.354998890613718, 
    -0.0845925650502092, -0.139971475950197, -0.232167210620895, 
    0.109502445644536, -0.184750303964564, 0.0738253740403221, 
    -0.336821402311247, -0.0533260335882523, -0.133298028068569, 
    -0.0888653522450377, 0.110401509019308, -0.0103510413089314, 
    0.0438782062110331, 0.0166907201641519, 0.0429131413321763, 
    -0.0316480159588989, 0.00249185117371743, -0.0674634577139927, 
    -0.064459170241587, 0.0470424118038234, 0.0838699744906719, 
    0.0680579411559338, 0.0836819667212148, 0.113844396229536, 
    0.126489856585399, 0.203679816070286, 0.109257580880939, 
    -0.0896948942358817, -0.00782749060577993, 0.475417349183682, 
    0.0970358199808735, 0.0633418468359539, -0.236354744891778, 
    0.423830368901519, 0.382196597187372, 0.179987700951079, 
    0.149253542806262, -0.14016092514454, 0.567021283789795, 
    0.276797808257161, 0.0698187984302458, 0.235561289130385, 
    0.483157297169895, -0.144185907436743, 0.320391266076641, 
    0.597241649676064, 0.140142129534027, 0.150651224787251, 
    0.0990071041280047, -0.33124769076417, -0.270825386804873, 
    -0.170126636140353, -0.238362445914237, -0.102224469131679, 
    -0.226648181260014, 0.0925775146944822, -0.241640698192595, 
    0.148882641194775, -0.20075670447045, 0.122446022562343, 
    -0.000172148003794462, 0.0541226831548792, 0.0108568849418425, 
    0.0397347845171197, 0.0300237320140165, 0.0564396005960385, 
    0.0455451346045715, 0.042909821912326, -0.0535612578243415, 
    0.0286848561764562, 0.0712634053240406, 0.0835153353902648, 
    0.131720748762005, 0.159576869220846, 0.106360950356444, 
    0.109304882325198, 0.232712334042496, 0.161869953676416, 
    0.0471469701113281, -0.00519142328752872, -0.124244639088096, 
    0.314029243629109, 0.576441922525873, 0.135789547427187, 
    -0.305150059936343, 0.291289300358905, 0.405134117285225, 
    -0.244351047840245, 0.0207527027868887, -0.174706554879632, 
    0.595516646627182, 0.0728131801278966, -0.0936092181077427, 
    0.214310843049677, 0.600449611729615, -0.0195255009505144, 
    0.539613794058278, 0.483676568969259, -0.253880739482398, 
    -0.213374900989241, -0.0476209973603929, 0.0814686240243575, 
    0.00954844364077058, 0.033016412095313, 0.0418010527943874, 
    -0.0641423672590742, 0.218065455531655, 0.000230003566050518, 
    -0.0674239344456788, 0.00113666669114516, -0.149907843174076, 
    0.0442186680613956, -0.0400351898211708, 0.0475156682930966, 
    -0.0973273274084001, 0.0143512603333906, 0.0263363246770813, 
    0.119983556380047, -0.11679256915466, 0.116888208586431, 
    0.0320680872260906, 0.206894276304796, 0.390564268017173, 
    0.000212395862811965, -0.0628222591722272, 0.0484311270208699, 
    0.240351022182796, -0.00721823971891569, -0.0988155189560264, 
    0.528198649879551, 0.432460550674245, 0.445134851251961, 
    0.452522549114487, -0.153001730010857, 0.627353565437459, 
    0.650377907585697, 0.584481076009833, 1.18409344332597, 
    0.404693641625688, -0.0955490919531027, -0.225371928590368, 
    0.288822858867478, 0.0404602087547513, -0.0240056371534686, 
    0.0494763149381804, 0.0709367306632786, -0.146504495818062, 
    0.0156501495241885, 0.0519549568922716, -0.0285788825935563, 
    -0.00498798534152405, -0.0662192896472751, -0.0101985052100881, 
    -0.0587866410054642, -0.0821007353133445, -0.0342780578482938, 
    -0.0190916036183746, -0.111318255202439, -0.060127684351162, 
    0.0160262814872383, 0.0293196805933139, 0.0381660887119721, 
    0.0283079127740162, 0.0503335724399283, 0.0247185287246568, 
    0.0236840343981085, 0.102604762925591, 0.12938947249379, 
    -0.104366270948311, 0.146218468338864, 0.271169750581465, 
    0.05458252574993, 0.169251815846204, 0.437761227835163, 
    0.147877187644767, -0.0145673953628661, -0.048170271589571, 
    0.380658453782426, 0.330656416849811, 0.143690534306738, 
    0.287713858571364, 0.551832789361811, 0.206585748022181, 
    0.0329741217686165, -0.0317601628652679, 1.22392965466169, 
    0.201450649908731, -0.148512315122697, 0.0812438577585156,
  0.508630892265, 0.196658117668859, -0.104426309473056, 0.200547127702396, 
    0.466504842680269, 0.11155333530346, -0.130600195973878, 
    0.142069551347206, 0.376896229979675, 0.0763960773295591, 
    -0.0840636320587171, 0.0195135936676615, 0.0589008275502836, 
    0.032697994736559, 0.00644315420496738, -0.0309977611006698, 
    0.031406507310321, 0.00448563726613302, -0.147471514441291, 
    -0.124027407129793, -0.196218324965797, -0.0208159718568814, 
    -0.160340229860541, -0.136657000523351, 0.130434092722318, 
    -0.206378996021893, 0.0357747063157244, -0.107154782882495, 
    -4.71609297289788e-05, -0.191644338651109, -0.0138460082946167, 
    0.0479728056902428, 0.0731631871619462, 0.131029125292298, 
    0.150812841415241, 0.101591502554297, 0.116179402749969, 
    0.217081202202549, 0.132365940637103, -0.0366659807087644, 
    0.348248902383499, 0.301115659972751, -0.0209294890200509, 
    0.122801755128836, 0.58247197710287, 0.366266457014407, 
    0.126350024300675, -0.27603405751519, 0.148139356168622, 
    0.615643946137231, 0.170515622698363, 0.0408379594185502, 
    -0.00425702668508696, -0.032196276818836, -0.186119412730934, 
    0.585067460531579, 0.407803190179997, 0.074806009378238, 
    -0.161019990084965, 0.131441252627812, 0.252659588093829, 
    0.0481171140305748, -0.0995529596005532, -0.122499540941045, 
    -0.103847004758864, -0.0199598351964321, -0.192316091822585, 
    -0.0426535189915908, -0.130115434611911, -0.101772873368158, 
    -0.130125978687292, 0.0132980585984297, -0.078045807889456, 
    -0.0276636644303908, 0.0109653363524891, 0.0658023709727634, 
    -0.126425359372248, 0.0777367137927279, -0.241394194019577, 
    -0.104232391967213, -0.0201010030979335, 0.0143837606835766, 
    0.0272475743185495, 0.044049937647347, 0.0647362922167152, 
    0.0458208144854426, 0.0163407991353414, 0.0475171433312666, 
    0.0243314405823242, 0.154663314786945, 0.262887959488963, 
    -0.0878711996395312, -0.135376674640339, 0.601739451832896, 
    0.286053050102638, 0.0369152256974845, 0.101209114188374, 
    0.149331187166846, 0.483166197141598, 0.536119644596736, 
    0.00468256088513927, -0.215115042556467, -0.27881872490433, 
    0.457134250326536, 0.594150086096953, 0.230160383102829, 
    0.364288538206253, 0.746857831752102, 0.080475980690672, 
    -0.0233269290522755, -0.278106113259585, 0.0861855675692025, 
    -0.311711046181279, -0.118158029847478, -0.284183084716578, 
    -0.257644523169363, 0.0429959270188118, -0.0152670000562018, 
    0.20246461375142, -0.22253404238565, 0.0170155781315245, 
    0.144726467847689, 0.141756418286698, 0.323252844910234, 
    0.473677676991844, 0.215719499197442, -0.0826223489369146, 
    0.171923370473821, 0.560125808947899, 0.23322169933602, 
    0.0566265717878818, 0.072741928355947, 0.0652176105737718, 
    0.127782081709281, 0.102542234977789, 0.0458007072297111, 
    0.0750914819211481, 0.0772400953785033, 0.114195438144844, 
    0.123495673921243, 0.0482079098201621, -0.00621776543596828, 
    0.0435609946151302, -0.0176035066726882, 0.0218274691174876, 
    -0.00646966257553785, -0.00955582929110065, 0.0570733449612991, 
    0.0769554457063877, -0.0356979196850954, -0.035551447940547, 
    0.0458985877653722, 0.263107846973037, 0.269241171052546, 
    0.192853561713557, 0.115039956784394, -0.11165266155723, 
    0.243613494282848, 0.35144227177435, -0.0940727145860577, 
    0.297305713027966, 0.94527943208252, 0.0372765726406099, 
    0.0345661305230764, -0.107743997190261, 0.681471329740631, 
    0.334364488056834, 0.210872442710802, -0.183841942488122, 
    0.606374493762304, 0.385167967032732, 0.299790870053201, 
    0.223883550180401, 0.0095578872587818, 0.268009219279845, 
    0.16908252183077, 0.160792288426279, 0.254497270407267, 
    -0.0771595537489706, -0.0851520383288461, -0.168282730456002, 
    -0.0203911454115577, -0.122519806676216, -0.0336835588782473, 
    -0.236185655046498, -0.0561557440830868, -0.224857236578551, 
    -0.0783275784823071, -0.214142082683894, -0.0714756704216714, 
    -0.0948734663507121, -0.0238400806578515, -0.0499759871822925, 
    -0.0722124571866451, 0.0540732795046411, -0.077096659262912, 
    0.0600422234944504, -0.131179536944681, 0.00394263215792612, 
    -0.0904501435699854, -0.0522110899953683, -0.0578861756573145, 
    -0.0576446012510125, 0.0277989686007563, -0.0275878718712172, 
    0.0330092791294145, -0.0940525818380872, -0.0194626079467129, 
    0.0807828500124043, -0.0737853468118168, 0.042540148624851, 
    -0.1715796396269, -0.0291015302190872, -0.121886928718665, 
    -0.0692380611252563, -0.0806198373421265, -0.0811640012100731, 
    -0.0340459103239085, 0.00213042121016091, -0.230463123394273, 
    0.103116836299455, 0.298789744856979, -0.211915160545758, 
    0.101825862506389, 0.574012625014141, -0.0319958808853483, 
    -0.231804093095335, 0.244911219419628, 0.298311723904744, 
    0.0108923017279395, -0.478802684961596, 0.421903537808622, 
    0.460559522893662, 0.091919542981845, -0.054272164896649, 
    0.138004850255174, 0.538131454097613, -0.0678138021724604, 
    -0.1174910006105, 0.447362716559078, -0.145271605193285, 
    0.0119176390130064, -0.372013377710244, 0.111524317321855, 
    -0.59543947559001, -0.278550183929273, -0.0741863528333015, 
    -0.199005084368861, -0.023440767541489, -0.409541178416859, 
    -0.079855948882094, 0.143285590842641, 0.148145587166523, 
    0.0634334917837849, 0.251711654497912, 0.446660168902408, 
    0.327319178958146, 0.192678955266173, 0.206071215693466, 
    0.343303174692263, 0.410327684710149, 0.362833884071031, 
    0.310370228270021, 0.308332838463522, 0.33855811988762, 
    0.330159258773373, 0.287717811505208, 0.28063314474647, 
    0.336912042499068, 0.356932412395431, 0.290630123129391, 
    0.27043160172635, 0.242171717346102, 0.183948713109544, 
    0.104190902288674, 0.0838070843542677, 0.373780540646732, 
    0.375025885001292, 0.102344977181922, -0.0299346036208389, 
    -0.130547970110126, 0.183953635336385, 0.489637311679305, 
    0.475913156838325, 0.16302143815915, -0.270015075287997, 
    0.0871394607817689, 0.403401457982716, 0.401904421142525, 
    0.326891871043744, -0.109224661807271, 0.534771494072175, 
    0.227720830207923, -0.0779001400092366, 0.269435418781186, 
    0.43672641233993, -0.0104832960389433, 0.501223528023026, 
    0.462721292320387, -0.253680522532059, -0.184601669395584, 
    -0.194452011718749, 0.395232980133458, 0.213328589380268, 
    0.161333616845265, -0.0740225539648369, 0.170219689179139, 
    0.230324405590338, 0.373943921722245, 0.14184507085431, 
    -0.191662661982897, -0.0773789727068815, -0.141339800880539, 
    -0.0188171068608559, 0.0378754340849868, -0.0650282271297668, 
    0.128696098235818, -0.0260919444109004, -0.0459909310314294, 
    -0.0586006545519041, -0.00684762998158837, -0.240209215933274, 
    0.0792305750364788, -0.0884867528350658, 0.0896373676793626, 
    -0.175413937404972, 0.101565274263049, -0.121853097431533, 
    0.0736204027384719, -0.25233627836031, 0.0043944272666753, 
    0.0404621474235117, 0.0322617555789754, 0.124066681948085, 
    0.191356059461195, 0.116708118572577, 0.064617319260808, 
    0.218046022672313, 0.205076583281357, 0.102068249386919, 0.1327804504784, 
    -0.211210260261881, 0.247477931494987, 0.669596326228856, 
    0.119566677898606, -0.0901548552004637, -0.0651920473705181, 
    0.552910128753022, 0.173953494519162, 0.30049592101802, 
    0.823217566606209, 0.270646716488345, 0.108103559381861, 
    -0.267228250065567, 0.167508943130009, 0.576882992504417, 
    0.220061345130602, 0.000724499361727527, -0.120832299098692, 
    0.179743972115451,
  -0.0367357716537779, -0.0756672282822745, 0.0155904273158738, 
    0.096208436842382, 0.0181278454811257, 0.0366968041926476, 
    0.138229134201456, 0.00629463763699478, -0.0428852442631418, 
    -0.106441647856774, -0.0200367791228641, -0.226192366252093, 
    0.0351690736793461, -0.208988160157894, -0.047265235003287, 
    -0.138492286416218, -0.0384327613201614, -0.0957459761207766, 
    0.0104093648415447, -0.227157436926268, -0.0165478870351686, 
    0.0562668721770693, 0.0527295169629686, 0.0723685580262644, 
    0.13171008847145, 0.116954494645945, 0.0900244472874486, 
    0.0865823973652526, -0.00232652258163857, 0.220559895147296, 
    0.406914620396718, 0.211826597749332, -0.153437490882035, 
    0.680942400033302, 0.207405228692987, -0.157775136741717, 
    0.310123096265009, 0.463799715956669, 0.0687875516785887, 
    -0.190516930182235, 0.528022704386011, 0.512140819735164, 
    0.237284015065878, 0.176161253916691, -0.34304683649717, 
    0.342588926305514, 0.337661951009921, 0.139670822347124, 
    0.635913753860911, 0.309339703540219, -0.0595928938141901, 
    -0.0125786325916286, -0.114965103888239, 0.0432177581108269, 
    0.223991782430962, 0.0748894181317244, -0.0029875572678502, 
    0.0210572929099798, 0.259946531006909, 0.00192401824504787, 
    0.00902796066815465, -0.0446902044684923, 0.0705898682929993, 
    0.0362047000907775, 0.0119892504551313, 0.00613458788152023, 
    -0.0351421463582836, -0.0204699426435271, 0.0567406149545707, 
    0.0421257622558344, 0.0364097953865705, 0.0481935936056699, 
    0.0282066459070448, 0.0429605567340183, -0.0113166027528207, 
    0.0258252446966345, -0.0327275071682309, -0.00964433360555679, 
    0.0440249735235078, -0.042230499445652, 0.0136165054148854, 
    0.15080142466606, 0.1819125937718, 0.0382174452459881, 0.150090589266496, 
    0.428201455795834, 0.176150855223279, -0.0437464978122819, 
    0.128971047615893, 0.386740875146356, 0.206052038620046, 
    0.103846640957972, 0.0765216135215721, 0.154607279403609, 
    0.164026628580462, 0.0941309691995703, 0.0610641149372561, 
    0.152783167060004, 0.158734964483531, 0.0679299723424651, 
    0.00582706731217193, 0.162687463923129, 0.255623558064979, 
    0.163065924426695, 0.0770621263788786, 0.000752685781018905, 
    0.252683264449493, 0.351795608059057, 0.148926239935377, 
    0.0459008646988503, 0.398053691104942, 0.177368260577686, 
    0.0034285358083017, 0.115972819721842, 0.339018902399939, 
    0.0454175952451026, -0.0616259453892809, 0.207342388452199, 
    0.066552281440636, -0.193834754049827, -0.153825778081156, 
    -0.277494504355621, -0.106775011737836, -0.0747761504195818, 
    0.0619056248365682, -0.291578955324126, 0.0452733983544926, 
    -0.0978635219712564, 0.0290657438937393, -0.271484696736911, 
    -0.037466378489682, 0.0939224451563082, 0.128334192912061, 
    0.0955086318199747, 0.081563493569148, 0.112378481245282, 
    0.124948459154271, 0.140886228412161, 0.121047083480412, 
    0.0410338419573309, 0.144603201040789, 0.259324353544802, 
    0.184803133127769, 0.123671611337213, 0.409028631885725, 
    0.318732697701789, 0.0844657799711163, 0.219981243968291, 
    0.50925211177938, 0.428191701537517, 0.175465191286058, 
    0.0844739061602979, -0.401579509863809, 0.779042623879396, 
    0.326460149883691, 0.0605684193906928, 0.0507881849290058, 
    -0.299036433995151, 0.190114269696694, 0.654658938645671, 
    0.593657441854137, 0.232103958025416, -0.27850454955898, 
    0.212176503149972, 0.472587160380569, 0.0818083469133572, 
    -0.229417888561908, 0.0387351482228233, 0.511461563187622, 
    0.520437117115763, 0.2956761392443, 0.120355900614989, 
    -0.242740269784876, 0.515956219169802, 0.425565005866791, 
    0.132524466779827, 0.306977844465089, 0.527305405729282, 
    -0.216827163462957, 0.0167312103900007, -0.371199817096371, 
    0.0973599204554173, 0.392207869161373, 0.334045036588536, 
    0.525296987301594, 0.416987036289181, -0.109716167885613, 
    0.25704128341411, 0.771947146888198, -0.18294915555756, 
    -0.121497105034817, -0.0628194458210428, 0.163197006925607, 
    -0.0347542604552622, -0.0381308852733818, -0.0132653664850393, 
    -0.0866309119551354, -0.0154681847405212, 0.00303234075351627, 
    -0.0261323792077543, 0.121136259094264, 0.0376079981823133, 
    0.133702493985029, 0.206190658538879, 0.106672859429081, 
    0.185678228485696, 0.319623301134546, 0.151851427401601, 
    0.102031453003838, -0.243593670537616, 0.331603355004168, 
    0.36903560349557, 0.121853500108941, 0.005048921740972, 
    -0.183253240352989, -0.0130283480035867, 0.517042617093564, 
    0.319531833318898, 0.237866859931975, 0.383052143621365, 
    0.0341997010597611, -0.0829601910314949, -0.097073019551105, 
    -0.0902874899297731, -0.0960302137262611, -0.0669640643410462, 
    -0.0906373614578215, -0.0204278433939228, -0.107115813401087, 
    0.0126256528957246, -0.0305755484031731, 0.0506013155675573, 
    -0.104476602633326, -0.0180005884527828, -0.00322054335545754, 
    0.0413525190768513, -0.0890874962309007, 0.0373302038406601, 
    -0.168857171134546, -0.0729315596600861, -0.00918428277618358, 
    0.0825995955936216, 0.131479315448692, 0.119658306914183, 
    0.0997457607927287, 0.0823756023570913, 0.153039828293561, 
    0.259177967343842, 0.200912932531841, 0.114565464807273, 
    0.110621066081955, 0.0470056148098726, 0.334120623708943, 
    0.465991070643907, 0.187003352598614, -0.176588148684118, 
    0.32354100165303, 0.634476245556636, 0.0741797800004068, 
    -0.235981569449853, 0.0812549108988871, 0.605435976301324, 
    0.103580581462575, -0.0544045816185171, -0.132143439315983, 
    0.286102695532049, 0.526644729923076, 0.267377750234335, 
    0.0326092531287562, 0.517151179797485, 0.292577978492968, 
    0.0788633441544808, -0.0350181912105437, 0.421252746032694, 
    0.243992570287441, 0.0186819064855498, 0.00836854436741248, 
    -0.336656203142277, 0.143195733251633, 0.363352870223076, 
    0.122375385947169, 0.0655762898719897, -0.0138718675537362, 
    -0.0363458632020508, 0.00954074413067706, -0.0337401992103667, 
    -0.115291193034022, -0.0264150242579353, 0.0409412868128911, 
    -0.101147679270201, -0.109991249447506, 0.0517546365841593, 
    -0.153029563785058, 0.0584223204776281, -0.273409985323722, 
    -0.0515040399651349, -0.101472323659491, -0.0932155330033732, 
    -0.0569053090380199, -0.163390147952543, 0.0122526361049579, 
    -0.038593910524981, 0.255226506657911, 0.160442552433035, 
    0.0142955067047146, -0.0805902015345941, 0.309405601186946, 
    0.329646555309375, 0.0966163163954484, -0.179809947631858, 
    0.123808142935105, 0.522097071130086, 0.208429438344031, 
    -0.22935397850089, 0.504562646866473, 0.702838320685436, 
    0.207425322622878, -0.0983794460411249, 0.35254944052696, 
    0.599002270193233, 0.255157820327872, 0.134062398115209, 
    0.841620419666241, 0.570143040190724, 0.362663401116982, 
    0.430171337414771, -0.555368576843291, 0.387918122095741, 
    0.661571854630431, 0.230159812305026, -0.268975244216122, 
    0.249386246512079, 0.204809976051195, -0.0486642120520252, 
    0.151864542240673, -0.219604099796482, 0.251125361724683, 
    0.14358953719968, 0.0388884249882226, 0.0542359554394758, 
    0.151298969983003, 0.0384184012474995, -0.0245703705904555, 
    -0.0269567867875684, -0.0270908624413934, -0.0248188794118058, 
    -0.0281771901520235, -0.00571925816732835, 0.0586398519591652, 
    -0.0597821379967515, 0.387260108278904, 0.0368082538845011, 
    -0.25624396104523, 0.0912154643265317, 0.791651996230635, 
    0.265957203498535, -0.0241981633037012, 0.0731712917177691, 
    0.853655186504904, 0.0592249767971393,
  0.000541992038743569, 0.0991037401321734, 0.0427192639353001, 
    0.0160711812567901, 0.214449071517264, 0.182371084315316, 
    0.0491415280713086, 0.158885299944568, 0.293252537650657, 
    0.135456210886983, 0.170921307723168, -0.185860684069254, 
    0.593584856059051, 0.316095460928353, -0.0409008819262922, 
    0.411474551212551, 0.39655564445653, 0.105208176002465, 
    0.697053336002791, 0.556325596729693, 0.287990143871828, 
    0.201816220366737, -0.226956229751156, -0.0123227068347804, 
    0.381018485150953, 0.390116717487978, 0.143219061907147, 
    -0.00614585029291623, -0.10332596698164, 0.135636048946709, 
    0.228109291047578, 0.281773614217301, 0.0750293361548641, 
    -0.040433316838301, -0.0189155678206515, -0.168721022636936, 
    0.00443236551860922, -0.0570086682420237, -0.0941641301224797, 
    -0.0639239654596657, -0.158086909003275, -0.0603763909397901, 
    -0.0559531799898431, -0.166182493516622, 0.133911694942633, 
    -0.0881685042891741, 0.0393423751089758, -0.0609666983777319, 
    0.0123730888724703, -0.153522667166671, -0.0388638159267198, 
    0.0701058081754365, 0.0696497910452419, 0.0711518423075443, 
    0.116728499635018, 0.0604977388627098, 0.19895841940918, 
    0.209839445625437, -0.0738270945785702, 0.0352843952917802, 
    0.562683727783855, 0.201969387262352, 0.23771154069272, 
    0.391045775157942, 0.619940280141984, 0.718091334603998, 
    0.224629722615403, -0.0616451569660008, 0.0771066772783001, 
    0.106200768339995, 0.0783581365870722, 1.01555286098994, 
    0.296652444758429, 0.0543508882696789, 0.156339145030044, 
    0.0346132269969094, 0.434200351020048, -0.129369821176217, 
    0.0193098637173694, 0.972652608562051, 0.234500323153844, 
    0.0249566896518967, 0.00112436877189337, 0.0120603161139762, 
    0.0256153269408892, 0.00536401966469312, 0.00777856903214692, 
    0.0841918340519442, -0.0252166797468604, 0.0760729286939012, 
    -0.165763930318167, 0.383466451766527, 0.180166870862464, 
    -0.0356745398293212, -0.164668181065974, 0.452725076947726, 
    0.38970900423625, 0.102969848722754, -0.0276535876269665, 
    -0.00589569862684547, -0.246106216342882, 0.623299097647754, 
    0.567150950977304, 0.254870683339311, -0.271170858224648, 
    0.628339052068628, 0.333011796214174, -0.0796679307462746, 
    0.47799537223591, 0.42296234220713, -0.116019796388572, 
    -0.0982762871801796, 0.0553847088734868, 0.0686363321003863, 
    -0.0112527890327933, -0.0288060380709863, -0.161879994698161, 
    0.00749850854159068, 0.0714016193149675, -0.144051454307215, 
    0.0216314310824319, -0.0447398899074698, 0.0304671309010929, 
    -0.109540234795778, -0.0173345915772643, -0.0782114167003232, 
    -0.0200731732119175, -0.086115311227356, 0.0647300518188695, 
    -0.0963936861319758, 0.0486810477095225, -0.0310177297780489, 
    0.0769216066007798, -0.0743919619435193, 0.0430354396303451, 
    -0.0518144714674296, 0.0267193837987703, -0.112203810151298, 
    -0.000914002692325166, -0.0342641113857012, 0.0385153151724674, 
    -0.0502199690486591, 0.0373165047461528, -0.0623275176642954, 
    0.00932650504088145, -0.0377660807626952, 0.0253219285787974, 
    -0.0511119119140431, 0.0275387322627167, -0.111394882575664, 
    -0.0152284569479231, 0.0195975664940338, 0.0234026422599121, 
    0.0167886268734681, 0.0297148831126294, 0.0354834708763017, 
    0.0385027474473487, -0.0625378672552408, 0.139981168804654, 
    0.127522155414758, 0.00940797772314267, 0.0705903624207916, 
    0.18760720345145, 0.178456437006323, 0.619641881321281, 
    0.419537968598183, 0.279568944468432, 0.279268726790855, 
    -0.144254025734921, 0.235675641992526, 0.686278121466732, 
    0.0114619750607998, -0.205512754437131, -0.353479751778757, 
    0.340135134609979, 0.653192814294339, 0.133978187783641, 
    -0.242391596508662, 0.032882352030923, 0.548999855857223, 
    -0.000178881795222432, -0.0307470975061917, -0.0973764197906256, 
    -0.151845057322419, -0.236564375030066, -0.157099008522137, 
    -0.10843228279792, -0.117650427256265, 0.0305027116019172, 
    -0.173961765148959, 0.0232926904481616, 0.0488793576852531, 
    0.0396815016162382, 0.0450280002618639, 0.0485950703482706, 
    0.0523702228075168, 0.0271328403849024, 0.122818678589453, 
    0.166917167324971, -0.210507813538722, 0.315943620615049, 
    0.321691290428892, -0.0444200134349135, -0.017515877169351, 
    0.453129398773742, 0.359387300895471, 0.385058213438812, 
    0.28664457952974, -0.16895438070569, 0.403822942079035, 
    0.352179557947232, -0.327115183696674, -0.00662040549374816, 
    -0.49559118165025, 0.669276916157997, 0.198814206640794, 
    0.0607973328880011, 0.386469501147038, 0.0922241669682823, 
    -0.182038920889205, -0.299149444597146, -0.0831790350393331, 
    -0.23411051364715, -0.214587288568219, 0.0524054748230525, 
    -0.137134562181845, 0.182127917131102, -0.144613445592951, 
    0.125495858714825, -0.250355094886054, 0.0312870462871043, 
    0.0867458441675002, 0.141065483073497, 0.247451338203463, 
    0.290080432836706, 0.28206150162158, 0.244701330664233, 
    0.217696386534662, 0.304420904727217, 0.351075360106803, 
    0.248811250173878, 0.188477300097408, 0.169356067531826, 
    0.162276864146975, 0.167165437856957, 0.176173166132466, 
    0.172840677925939, 0.164046513651692, 0.197315842724422, 
    0.191073650970399, 0.109122796749017, 0.0945604426169508, 
    0.0945882436830731, 0.0868333864790839, 0.0956180263998562, 
    0.0675765761605742, 0.0493326325869592, 0.122994320315902, 
    0.105530564952704, 0.0219917808042194, -0.0346382126850044, 
    0.240323688867027, 0.235419178587735, 0.150777264419667, 
    0.256605816474426, 0.141432487612513, 0.199593018083401, 
    0.593009629861698, 0.111527573249757, -0.0618130837623966, 
    -0.0774409263481173, -0.24150479015988, 0.788177038648332, 
    0.183498920940707, -0.14730211479359, -0.11538069257154, 
    0.742406239490553, 0.370063836895062, 0.105482350418973, 
    0.342447034565457, 0.285134130693703, -0.0804676836025739, 
    -0.17475935299508, -0.173031822313088, -0.0855514071468101, 
    -0.124431270268349, -0.0518187049880682, -0.014378782973703, 
    -0.0981573336589776, 0.0570496154814017, -0.154042064326502, 
    0.18052632906405, -0.035923863551483, 0.0935904523361529, 
    -0.181727230442431, -0.00741204689627355, -0.135046487362718, 
    -0.154220007816392, 0.207157824416934, -0.14772451934627, 
    0.0890998310010422, 0.0170270768977738, 0.0334186731233861, 
    0.00744494288768813, 0.0167360240217157, 0.0143749992283497, 
    0.0192617833401172, 0.0315243382766915, 0.0372703588367709, 
    -0.0440674243961831, 0.0610248717367241, 0.106143313524896, 
    0.120509020705089, 0.176497972323874, 0.176323638510116, 
    0.0828057635051548, 0.104250403538152, 0.377096473844532, 
    0.212621178746755, -0.0883578747351079, 0.458046786132941, 
    0.362243188997152, 0.0956758387562498, -0.212517358426317, 
    0.196327714251134, 0.595454662220516, 0.244994869937172, 
    -0.0915022507629237, 0.185657531412672, 0.401560109012885, 
    0.301757188225542, 0.224272347481611, -0.177676935580592, 
    0.338890678635574, 0.719765678955401, 0.118129630913279, 
    0.0308021141687709, -0.0724673677513516, 0.263140464898417, 
    0.429739111221198, -0.143832198785857, -0.0593577500592091, 
    -0.00397775670019054, -0.184317653091012, -0.064457207192416, 
    0.040931385663765, 0.0143892482744206, -0.00314165151838054, 
    -0.0967403343248487, -0.145620798184728, -0.175961234221161, 
    0.0226956450074638, -0.183472044766131, -0.00689026661944926, 
    -0.121626520791561, 0.00167328809416596, -0.280313787740184, 
    -0.0801644987175671, -0.137350135937285, -0.254708250538388,
  -0.136267101028481, -0.103941649461614, 0.630356781812512, 
    0.558187797103876, 0.297491779210931, -0.221385632794897, 
    0.139899125685712, 1.31130778236871, 0.121370651365175, 
    -0.0877354755344076, -0.182377697758961, -0.171583563347457, 
    -0.153044591781064, -0.178081683559778, -0.125036404727037, 
    -0.161819603917138, -0.075093230322525, -0.153711790356864, 
    0.0205073263238531, -0.210406403299771, 0.0754776006084081, 
    0.122772560689002, 0.095864037617989, 0.178658278919457, 
    0.222042143692917, 0.153499033279541, 0.202910266815705, 
    0.333225631310379, 0.172985936016426, 0.0226144136047851, 
    -0.056488021206803, 0.384646299523372, 0.336007318029583, 
    0.119274503423292, -0.111582660293934, 0.138760202260511, 
    0.434788641047687, 0.264452381280524, 0.114044241854375, 
    0.0193864454161937, 0.139080722682804, 0.367749587304325, 
    0.289635762680879, 0.15452981759611, 0.212382849026624, 
    0.414169542059502, 0.335377294281437, 0.138407928374834, 
    -0.0884456553858955, 0.342797935687593, 0.434285406682853, 
    0.104000907670707, -0.0236827824199935, -0.0452827743442717, 
    0.130540542071276, 0.353655697851147, 0.483959350583896, 
    0.267218695918659, 0.0837279803098705, 0.539897144819939, 
    0.283953012347265, 0.0747519611282973, 0.204412997848523, 
    0.268310740103051, 0.070132029868242, -0.252333031187077, 
    0.468066878097383, 0.143927054768777, 0.0552094102485887, 
    -0.0158595765810023, 0.0650233137966556, -0.23339437834011, 
    0.265776219652301, -0.217814246264514, 0.0288678172172064, 
    -0.240806130145353, -0.0540231878153962, -0.0991474858174997, 
    0.0479746364816194, -0.402056364097439, 0.00169136368628722, 
    0.0676849702377306, 0.0902962923897224, 0.134346347879944, 
    0.141684811688944, 0.0894721242225453, 0.110515855177864, 
    0.143775876949636, 0.121931637081962, 0.0517349016507827, 
    0.0909566082871543, 0.111263143724182, 0.100663838146865, 
    0.127984036349486, 0.167995436532353, 0.130514940018461, 
    0.119938992489703, 0.262892635484728, 0.175034411125551, 
    -0.0880002773603458, 0.261381210592198, 0.330932429864792, 
    0.0215698335145425, 0.408676667503103, 0.461201989398256, 
    0.110544710678018, -0.0445095197794332, 0.240942669054027, 
    0.387458495458144, 0.478105631234426, 0.387649688413833, 
    0.107214089482442, -0.0287689127252566, 0.0980482137363138, 
    0.562431948051919, -0.160893014546996, 0.0206985314720905, 
    0.827795392374523, 0.279222426664151, 0.0491635557533615, 
    -0.101266208359576, -0.228045219916934, 0.0965085626428098, 
    -0.117285866766185, 0.0219868244244864, -0.157810093203984, 
    -0.0257706087979187, -0.0655149328447671, 0.0220611031915836, 
    -0.216199655806136, -0.00944808296968708, 0.122093203950803, 
    0.140375546674327, 0.168514545952001, 0.285876798644959, 
    0.304150000685147, 0.230184780717491, 0.197645476141286, 
    0.228841983811383, 0.277496060715796, 0.322720413384072, 
    0.303078197542989, 0.272697337456065, 0.275397069098856, 
    0.299362513627574, 0.334288252647087, 0.311946433311882, 
    0.170959492563071, 0.115054579548703, 0.55174447599083, 
    0.321828791694005, 0.0437385464846431, -0.123674456332777, 
    0.437213283816897, 0.397547835741834, 0.192320605705152, 
    0.127565966194863, 0.16617196634268, -0.206787069715482, 
    0.647205192104881, 0.387845951440853, 0.129583421575527, 
    -0.266165609157805, 0.589713157736903, 0.283646100960918, 
    -0.0600187517549448, 0.210233229240323, 0.519979872349241, 
    0.210279134402522, 0.0205086186411167, -0.0910163100637293, 
    -0.151725595139066, 0.248866553052542, -0.0199641834565213, 
    0.156119886617383, -0.328882347827794, 0.0193774405322866, 
    -0.0661680983242371, 0.118804774344714, -0.284786010714833, 
    -0.0407423771320046, 0.199898566725231, 0.161367793592095, 
    0.104230736294074, 0.16102285919043, 0.308071947782538, 
    0.375666317171659, 0.323188708407597, 0.241631392414741, 
    0.223330631016687, 0.322838873285501, 0.371907492681706, 
    0.39021206612009, 0.456075876777483, 0.467699640380568, 
    0.387554437219305, 0.338178846136673, 0.353475972468805, 
    0.368612994635019, 0.376175415357678, 0.340325216510514, 
    0.333103080203753, 0.454138422562049, 0.45338392768361, 
    0.197818523163237, -0.0569235710817328, 0.307382961491133, 
    0.426490658969106, 0.465546649935371, 0.241405157685231, 
    -0.237423348022335, 0.067479677143462, 0.591415828511551, 
    0.143015511154181, -0.115025450074012, -0.0338237935906227, 
    0.44784598307092, 0.257782384800897, 0.264941379608307, 
    0.595633404446346, 0.173262381738397, 0.0260546373488675, 
    0.0696202765284292, 0.189590256323732, 0.20701871680574, 
    0.0812282912780334, 0.144635547958863, 0.388411574339335, 
    0.0613631085573731, -0.00928431804920629, -0.0621902140382945, 
    0.0414702001526823, -0.0830763638297934, -0.00199271833253475, 
    -0.080489141143057, -0.029897160819117, -0.0580650808498959, 
    0.072810109591962, 0.0817901497662025, -0.0947603861466783, 
    -0.19545065187314, 0.198061704389538, 0.414095994309294, 
    0.172143314388413, -0.118359778636043, 0.340395774805451, 
    0.399729763298219, -0.110154332828202, 0.0478481499533048, 
    0.104767388534774, -0.207131890304539, 0.749981394955813, 
    0.22854681781609, 0.00809053140147246, -0.0101151834107562, 
    0.330499971131467, -0.0269714711993305, 0.293160794844814, 
    0.905575101388854, 0.465892540147566, 0.164171755527938, 
    0.230919131074774, 0.128712591223582, 0.416389352033359, 
    0.425110299670508, 0.0881947781158187, 0.0168067487045662, 
    -0.0257825345103134, 0.132012526386742, 0.124656568670243, 
    0.0766678731753961, 0.0286804773701071, 0.162397726682401, 
    0.267624010534453, 0.0790360029110675, -0.0119103278110367, 
    -0.101421731276312, -0.00164335009723586, 0.163980669233916, 
    0.0297766857509894, -0.0298795223208618, 0.059009747627994, 
    -0.0221432439185048, 0.0337709919656821, -0.0280977342583407, 
    0.00984786515325428, -0.13404281597492, -0.0295093971244264, 
    -0.00848653009142238, -0.115256061557437, 0.0475251140986401, 
    0.126470622832729, 0.047460473318112, 0.0819095400863698, 
    0.331778023281172, 0.166572766783819, -0.0155278064862535, 
    0.0591182218206247, 0.406384377043154, 0.125714266437156, 
    0.0977069992234652, -0.170244125008997, -0.0523458175839268, 
    0.647466416156577, 0.360343221421976, -0.0314102327809462, 
    0.40052425563357, 0.511956966428634, 0.318236525580056, 0.18522743843251, 
    -0.0139483168891189, 0.272491476932731, 0.00329471110848838, 
    0.326638534388639, 0.728442040670228, 0.254933019522038, 
    0.113019275662774, -0.0673899142741561, 0.508109561683657, 
    0.0507542416372549, -0.158773264501154, -0.177086834532854, 
    -0.0610341375772002, -0.164142935659907, -0.226162138566694, 
    0.0559344481165786, -0.135315239191268, 0.0107038012543152, 
    -0.27052059352401, -0.0520415065673615, -0.154890833586841, 
    -0.0910705270285937, 0.100139978845354, -0.125048652999938, 
    0.0770137190940342, -0.0465454809619352, 0.0216234030491489, 
    -0.06106377378505, 0.0238938406533917, -0.173352286626168, 
    -0.0117381588876267, 0.0230685650392498, 0.0400644581058027, 
    0.0776815776432172, 0.101491844553976, 0.0640038045208082, 
    0.0308398738721519, 0.0628091002066828, 0.0365647916346686, 
    0.0551068798065143, 0.338813954836927, 0.150412374591578, 
    -0.0548827504390669, 0.0935733393392005, 0.00255799028352878, 
    0.685771849391062, 0.460002346491179, 0.118785104223894, 
    0.759687662806033, 0.272842009570545,
  -0.0222084365384191, 0.0590261308377138, 0.225294998429803, 
    0.202703233024382, 0.158050996353567, 0.153523186720456, 
    0.267868190857024, 0.346630639018122, 0.216222890628815, 
    0.104203958813693, 0.0798748064736721, 0.0650419208618599, 
    0.0734014416597312, 0.0655414188114597, 0.0701033441109019, 
    0.0613130467910747, 0.0697845998226349, 0.0643254612671665, 
    0.0777942982770491, 0.0224845814704663, 0.190547777000005, 
    0.175283548121201, 0.342317075932483, 0.206398894479174, 
    -0.108699783535861, 0.0906451815638774, 0.670183269495696, 
    0.0651759511846562, -0.247608808554932, 0.158255883793615, 
    0.470736790589624, 0.0566807005575724, -0.0137411778418219, 
    -0.133299322627465, 0.234219298542721, 0.121895627480083, 
    0.397401550540514, 0.892305813854, 0.465600139006513, 0.115873540748669, 
    -0.00646437231129803, 0.0909283148856103, -0.295948036718292, 
    -0.169096511106999, 0.413624171855815, 0.225065094138834, 
    0.115929089133217, 0.41323023559395, 0.350821406177964, 0.12771691249173, 
    -0.0767647643204768, 0.301209987952383, 0.268021786694612, 
    0.00875240895337506, 0.406215401498813, 0.441103515692037, 
    0.13364807393613, -0.0548351725525326, 0.550084496477272, 
    0.297936092250787, 0.0840928315612907, 0.00485229426946168, 
    -0.311115230456389, 0.414282897002795, 0.616016999841758, 
    0.236957101181103, -0.264838535253704, 0.0776906437343475, 
    0.417815490489841, 0.0763343734853093, -0.0609972527179325, 
    0.12603156913442, -0.514814905748132, -0.0629750941764016, 
    -0.116759447919491, -0.332888629962565, 0.156847448312755, 
    -0.035633184002393, 0.225505544117641, -0.226565645684317, 
    0.128533525051087, 0.0728447363420771, 0.0847309676413006, 
    0.171181640475554, 0.192888983590482, 0.121067174030158, 
    0.101726865171202, 0.118142257351966, 0.15472318176457, 0.13794052066335, 
    0.109586065437426, 0.0702359246589426, 0.0770911599811103, 
    0.103136315429603, 0.0827812416000215, 0.0824937890133354, 
    0.0395666951996221, 0.163444783627715, 0.3137463416357, 
    -0.182431940508973, 0.42450487487608, -0.00220115578240344, 
    0.432638563924975, 1.05736575432311, 0.395876776320361, 
    0.0267289932247399, 0.295534247109377, 0.809361440645957, 
    0.125950868160396, 0.021444534594444, -0.310492877340946, 
    0.395444894562847, 0.55285412299709, 0.174869891773404, 
    0.021779496877871, 0.0402478665652722, 0.125149114381923, 
    0.387854904446349, 0.0633696622262822, -0.130293008596391, 
    -0.165322497762595, -0.0708281867670541, -0.101424348151759, 
    -0.107010106753811, -0.0885834758899139, -0.0700325074421317, 
    -0.0756878387696728, -0.0145968019483316, 0.274668059956982, 
    -0.0944571271195611, 0.370326629918134, 0.31248403730341, 
    0.0692954265969538, -0.24620620768926, 0.041969941700476, 
    0.498323961853851, 0.176107162286339, 0.0968807264295473, 
    -0.235028860918091, 0.222403025620047, 0.376084715574543, 
    0.196583960904485, 0.111586264602103, -0.138090962179809, 
    0.285352762547409, 0.263964367543439, 0.0636790636185111, 
    0.163143460326792, 0.390334721679508, 0.0947785347860217, 
    -0.0483291526230007, -0.0346986954689629, 0.00676211512573856, 
    -0.0248929476794934, 0.00312372445548806, -0.0322400573413273, 
    0.00018996585528587, -0.00067752590424186, 0.046333325545748, 
    -0.080062549382645, 0.0749900716484373, 0.146315306703953, 
    0.0661982764574651, 0.252407844065402, 0.232436067894829, 
    0.0464215008425304, 0.164693193905454, 0.354096993245578, 
    0.27027119528988, 0.0837726412921471, -0.0505980126248004, 
    -0.287182828238929, 0.275612983091746, 0.652366458208373, 
    0.130517890377741, -0.118688202681536, -0.0878989777000191, 
    0.297707602198211, 0.535931959658302, 0.313171843878758, 
    0.0194696638622261, 0.0620548534556022, 0.240732782514162, 
    0.0313304836278848, -0.0613646185082007, 0.0703141652194592, 
    0.150111607691552, -0.146306516264822, 0.0746015431728807, 
    0.0443278134855353, -0.177227914959523, -0.0633157308907322, 
    -0.102996858253292, 0.0231602223499337, -0.310457357680355, 
    -0.0237578629802277, -0.0861958164031937, -0.193356480824714, 
    0.185797837010263, -0.239492966689701, -0.00015375091911915, 
    0.0470690991001913, 0.0586888865441082, 0.139387553701697, 
    0.185498783322757, 0.126037061598077, 0.0836208749109648, 
    0.109234962412607, 0.158282089301636, 0.38932705158691, 
    0.259296104007067, -0.0939872262804238, 0.0983693918886733, 
    0.663490063194536, -0.0126125472047114, -0.0737218984701686, 
    -0.142962255278218, 0.563433104787149, 0.273459454300237, 
    0.117907374884439, -0.1615252151008, 0.01518120699566, 0.356028567012019, 
    0.498751319273132, 0.138860147495934, -0.150303601797852, 
    -0.0349407417593657, 0.301905248747044, 0.290041909132402, 
    0.374369327250375, 0.189112218269352, -0.0556650086935906, 
    -0.088108875709764, 0.0517942768309551, -0.148917704541683, 
    0.0313364102051639, -0.0162100702252904, 0.102577463442849, 
    -0.0397684032976028, -0.099638380393034, -0.140706417787136, 
    0.0720763124411207, -0.143874181411472, 0.0491777885254838, 
    -0.14149798874044, -0.00886532381975159, -0.317423364413333, 
    -0.115186928010827, -0.000935315219612973, -0.237801484495324, 
    -0.0229862219658486, 0.0919971206412724, 0.0097823363066866, 
    0.0585451980912166, 0.261018485339848, 0.0816400054464401, 
    -0.039540191544303, -0.0466135682677501, 0.0666546446690569, 
    0.405661715704761, 0.311829749024944, -0.0973396019099789, 
    -0.096721445758722, 0.454782670365724, 0.577196896084373, 
    0.233473272372027, -0.270628440829116, 0.217413019943006, 
    0.565934270545574, 0.0971888848213063, -0.0637096064288088, 
    -0.244876855683751, 0.177435679953133, 0.422509040941992, 
    0.00639001010497081, -0.271817901896381, -0.042296076783247, 
    0.522991340286564, 0.0881978079535969, 0.0836009463545851, 
    -0.303166097982148, 0.0589970417648792, -0.319957642134396, 
    -0.000594968562841455, -0.302950777711872, -0.0210000490652912, 
    -0.249742057932808, 0.0352304433476775, -0.270545134844897, 
    -0.046625874207143, 0.00527871449143226, 0.0319817619564861, 
    -0.118853558424378, -0.0642446173825825, 0.0862038142258117, 
    -0.0585325689699926, 0.0309918430232931, 0.0565042039423851, 
    0.0629373982563961, -0.0502004002854303, 0.0164738370105631, 
    0.0741557878529832, 0.094273466273365, 0.0750410985994854, 
    0.0703956382064728, 0.0815219238199683, 0.0872414793695539, 
    0.0739451886646646, 0.0741882384212728, 0.0862261820961494, 
    0.101899909652616, 0.0850275270747374, 0.0860622633889277, 
    0.0946957840955793, 0.101150143709392, 0.0865049683235222, 
    0.0910159199774215, 0.111837381842856, 0.103003822082636, 
    0.0627424779463968, 0.104719066764595, 0.127453452875879, 
    0.123766156872917, 0.162997959715935, 0.199402121738402, 
    0.15455238362181, 0.146873236056476, 0.197182903559813, 
    0.114234303056286, 0.0700456572236123, 0.458418024160379, 
    0.288562767555515, -0.0338243502142762, 0.437300164038821, 
    0.366803185353341, 0.0788601095752938, 0.209355470029569, 
    0.479467128398098, 0.325644885192001, 0.239255382822267, 
    -0.044234799904686, 0.640279795211076, 0.00169536368897774, 
    -0.165249505685456, -0.0219368620663981, -0.204235902490296, 
    0.231081911610981, 0.211235353600865, 0.109983160503897, 
    -0.168112782616482, -0.305143835826014, -0.387582788697315, 
    -0.0730719255549102, -0.488047887980692, -0.169629936310488, 
    -0.20911111709071, -0.199742325638689, -0.10680010958493, 
    -0.0635406434148395, -0.477794493543168,
  0.141429341392302, 0.157438667273824, 0.1155234413055, 0.152584719379137, 
    0.0731492571220486, 0.169144300127134, 0.365057627865474, 
    0.135669428324306, -0.0337584835984572, 0.00201161870669247, 
    0.507641147444863, 0.221104039617576, -0.0951655390327113, 
    0.49420397220745, 0.31293148047655, -0.175188319866496, 
    0.363546987715977, -0.375158194812453, 0.683759281995973, 
    0.0913944103658632, -0.100063476761748, -0.175960986895621, 
    0.0963689029851834, -0.00104189021570761, 0.12208301499144, 
    -0.0486714957351876, 0.164477367266791, -0.208335672635023, 
    0.0926028482879096, -0.195328774518895, 0.0064004557712966, 
    0.084445109826633, 0.143372748341258, 0.155182310159412, 
    0.12380353517273, 0.143742404584311, 0.0935293578404298, 
    0.107319506554251, 0.232567663286718, 0.145896394129469, 
    0.110222159881008, 0.124689692656526, 0.126154141933044, 
    0.121426708939083, 0.136907594294641, 0.136289609017534, 
    0.145173484926096, 0.162169008766008, 0.139926880680614, 
    0.115236339273474, 0.145579187934442, 0.157612252987878, 
    0.135071889953342, 0.13951908533065, 0.208382394607264, 
    0.179203189073784, 0.0790101290940818, 0.052683621366823, 
    0.224675081463191, 0.207443302623724, 0.26190375476964, 
    0.171214285840721, -0.0744182389451059, 0.012954403438906, 
    0.743470482057892, 0.160704705783745, 0.0779295911235082, 
    -0.369708350901911, 0.22395924733513, 0.542769521379103, 
    0.317007297933223, 0.365775125397548, 0.291571749317152, 
    -0.311860556429759, 0.226272432560127, 0.426533917695487, 
    4.5564570851947e-05, -0.408895579627564, 0.394978381150087, 
    0.81104910555662, 0.348521255295474, 0.113571504479989, 
    -0.0310335723859027, 0.00853079568373969, -0.0997257487291201, 
    0.0227596576031649, 0.0594484828897039, -0.0361657248058027, 
    -0.0566672870603182, -0.124401503182736, 0.185948896148264, 
    0.137700085003523, 0.0167170574659874, 0.127123020274243, 
    0.214150352649763, 0.145571146333219, 0.132414973393565, 
    0.172781647794435, 0.201992796827207, 0.240621564259421, 
    0.15461955644385, 0.0301043040074443, 0.0483740138429539, 
    0.295471884291503, 0.216439615213693, 0.0892884797039317, 
    0.0563333189495952, 0.219818996415422, 0.162509474082798, 
    0.0434239739146929, -0.0608660904748168, 0.00700871959247579, 
    -0.0120441060835113, 0.0148996888833747, -0.0521384684012359, 
    0.000472248516537752, -0.0198716750516273, -0.0356765702808659, 
    0.10273898751593, -0.0600364433681093, 0.0824917044167065, 
    0.149535209152618, 0.0587861669144889, 0.0850197967311997, 
    0.206463558089627, 0.122148896464994, 0.229532070984358, 
    0.30357500422232, 0.0739349112208863, 0.0537901689156066, 
    -0.0695828932959101, 0.770210730893267, 0.10994777028384, 
    -0.571264127577697, 0.150235261418423, 0.648635314222024, 
    0.248196153595799, 0.346273872461841, 0.732416573125848, 
    0.312153535833542, 0.0284448088343253, 0.332503247024468, 
    0.225888938101379, 0.192759883429906, 0.148893265475584, 
    -0.149660956134131, -0.286050845215174, 0.0160391083336793, 
    -0.22531815171594, -0.0578691057824664, 0.0270914233027819, 
    -0.316048168520212, 0.329537936358322, -0.183222205200837, 
    0.0552949490551833, -0.145479585290527, 0.0169311142384827, 
    -0.07783780673205, 0.0923284958093362, -0.244596310404794, 
    0.0679470282379505, 0.064617795419829, 0.0706439508616553, 
    0.0552512281859177, 0.0621992892130421, 0.0649671565871896, 
    0.0680039927227844, 0.0277414051114671, 0.0507563367644509, 
    0.0232832243573824, 0.0345418621065624, 0.0937242959755268, 
    0.179122667713182, 0.149215493164799, 0.0830368515176679, 
    0.0496366013871767, 0.16184721395855, 0.218982827589168, 
    0.280455372467159, 0.272311024113069, -0.250414308181563, 
    0.560636647089793, 0.392349525983455, -0.0666153876192995, 
    0.566472475598897, 0.375352317552471, -0.0375392093301104, 
    -0.37101238438682, 0.786154966073648, 0.328998019176316, 
    0.0399150902424155, 0.049852936915206, 0.0556574224457654, 
    0.044216056401589, 0.0545023027565595, 0.0499421110679054, 
    0.0498338629435059, 0.0664338397006035, 0.0414589890146301, 
    0.0283519937080275, 0.0791485444119671, 0.0910978815346252, 
    0.112844872042571, 0.15440089053902, 0.172588044944007, 0.14989080001599, 
    0.135964555351277, 0.171052248748286, 0.169970218216707, 
    0.145056861401264, 0.185834742897586, 0.185852152587478, 
    0.162742180517985, 0.149811905416663, 0.201802602951849, 
    0.278129226374746, 0.182072578183969, -0.075845746764357, 
    0.550901486312743, 0.219031771146509, -0.239896632572215, 
    0.229039405878231, 0.637157059470486, -0.182222958997276, 
    -0.100566147469157, -0.46377709406489, 0.525074169020962, 
    0.632376438914994, 0.268918530397818, 0.0941815799601124, 
    -0.0628271647962438, 0.225623838646756, 0.0446430641392749, 
    -0.112079142143052, 0.177717294654587, 0.166169842836138, 
    0.19663298987445, 0.219623836511423, -0.0455212622168009, 
    -0.111661359766848, -0.0959336810404967, -0.0697716359161122, 
    -0.0822338665401064, -0.0873007401492804, -0.0628246330015938, 
    -0.0886686887723133, -0.0258957363187976, -0.0835421379386205, 
    0.03723326036033, -0.118326502261575, 0.0730020289215319, 
    0.125947165624442, -0.0137982748466723, 0.19233356980535, 
    0.23577337476864, 0.0700408154820736, 0.00423541441267855, 
    0.308117298692726, 0.149208670210015, 0.0446833647084067, 
    0.27943432975426, 0.216958987319604, -0.250735880592351, 
    0.109705621248799, 1.12720710148565, 0.114093928139309, 
    0.103210158664468, -0.443961207854149, 0.249578480823376, 
    0.190818029456867, -0.417862474318906, -0.104651588886667, 
    0.0643418063035609, -0.156554431062343, 0.237458040758686, 
    0.232654167517427, -0.0518690047357464, 0.327231209084431, 
    0.134597234497282, -0.175617547429765, -0.0655509197529703, 
    -0.139150756689092, -0.0365609568087906, -0.145835390477029, 
    -0.0842555774979406, -0.135853495074795, -0.0973836103811583, 
    -0.0945385201561136, -0.105785668584307, -0.0984697073935889, 
    -0.00465042073346106, 0.151942642595917, 0.157445107133435, 
    -0.0346447425279368, 0.268057127926501, 0.416150201786518, 
    0.147912301646672, -0.0496573826425822, 0.301099015128922, 
    0.314904370528387, 0.122717608642725, 0.079728983675292, 
    0.10851742236733, 0.133622953785638, 0.115834411048855, 
    0.070088892755581, 0.081804627164674, 0.124467844589301, 
    0.125428690125558, 0.0586387102482287, 0.0419686081347421, 
    0.161485893458221, 0.185139740020312, 0.152381357468639, 
    0.316944201441132, 0.230398012607038, -0.0672505764687245, 
    0.299415003530353, 0.442073153582679, 0.00126163458439077, 
    0.0497952646266338, -0.147324351264704, -0.0351399643979709, 
    0.376050872513588, 0.675215909965111, 0.146251929166931, 
    -0.104273968486968, -0.0376791004121163, 0.584567164320385, 
    0.0159067264495097, -0.114337234737839, -0.0801743053637186, 
    0.269983176982352, 0.0839021791817493, 0.0744030454762011, 
    -0.1650557344836, 0.158579047697523, 0.220875442058868, 
    0.0559698322567761, 0.227380618264733, -0.0934678442189786, 
    0.174728935702375, -0.305497870413154, 0.0339323891712222, 
    -0.291149371654835, -0.115856675247855, -0.113107133011822, 
    -0.183602129427984, 0.0929340062023203, -0.229512454513315, 
    0.0448211432943312, 0.0456500262681498, 0.067548395338366, 
    0.0293252306250027, 0.0499504290009302, 0.0176314106625621, 
    0.0179738005246989, 0.0655188915954909, 0.0878398754372816, 
    -0.0114354030722308,
  0.202148209217407, -0.0368867370833201, 0.143295568476279, 
    0.196541644187939, 0.000563827520277949, 0.0246066050967842, 
    -0.207354872584953, -0.0145551519543404, 0.205118886451911, 
    0.195335975210859, 0.214797120655923, -0.0796153940556142, 
    0.797078870753675, 0.520434334981229, -0.0114272913935138, 
    -0.084240962034184, -0.401666412041243, 0.806396784098073, 
    0.1815716892053, -0.112234786523673, 0.0572417548050205, 
    0.425826358599368, 0.180341480932798, 0.72525048370028, 
    0.632390958517696, -0.0845315268844462, -0.0419851944291486, 
    -0.439670583892029, 0.125517083385348, 0.741876205338295, 
    0.295249151264677, 0.0771886999072208, 0.592901098541295, 
    0.299405838078865, -0.212397049620738, 0.272421726918823, 
    -0.412999928381505, 0.120086927590396, 0.313470935691573, 
    0.0894149099072524, -0.0303738297857766, -0.0209284072560708, 
    -0.201546550499026, -0.144638977923431, -0.042792578785505, 
    -0.162766757222022, -0.0531870278002468, -0.0697002955260972, 
    -0.0764515134429065, -0.0805511687949629, 0.0978235979090789, 
    0.0438554111621529, 0.0250646046405203, 0.138399611044888, 
    0.10961866909006, 0.10311653195214, 0.0871475649301593, 
    0.0409161898435067, 0.0363966365160111, 0.0469108553417596, 
    0.091793926815234, 0.116162482752326, 0.106332632421442, 
    0.101565395906936, 0.115544036093596, 0.105309515611769, 
    0.0846324290116346, 0.103147256565291, 0.117219738581979, 
    0.100662029988389, 0.0577278275566787, 0.0487613912065658, 
    0.068398194187998, 0.0726287728991654, 0.083861005856454, 
    0.0489530649019081, 0.0210013315722337, 0.111280178590583, 
    0.101180305068246, 0.0424954762645536, 0.159763204436562, 
    0.0433202755046288, -0.0153364081292813, 0.0979739751500946, 
    0.432453942199965, 0.437453458697094, 0.0897783192461242, 
    -0.0964523254918819, 0.0343880586866719, -0.187559477442497, 
    0.148804181419826, 1.0863632031692, -0.105134889632016, 
    -0.213571427172579, -0.326578830726029, 0.900555378385435, 
    0.210287421560639, -0.0737135469506338, 0.613965537847977, 
    0.0246927248946145, -0.36804330030811, -0.157974536003288, 
    -0.0270557482105241, 0.0431772836370159, 0.0097833513978345, 
    0.124271403184409, -0.106224634807459, 0.0804316359288838, 
    -0.193213535782126, -0.233443329312965, 0.0261366085836916, 
    -0.121102835738344, 0.0555423638719345, -0.137630469768867, 
    -0.0151988866126736, -0.14047456135787, -0.103466845439221, 
    -0.0276020909786265, -0.111611472075343, -0.0170145235986686, 
    -0.00860578179678282, 0.0297527000562432, 0.00553978889180175, 
    0.0192804090521572, 0.00724539611162956, 0.0152156916617442, 
    0.0112960994541422, 0.00237590911184823, 0.0418054851868365, 
    0.0483840857702109, 0.0235370253398697, -0.0534467273520396, 
    0.012741395618725, -0.0178596447893002, 0.0176948748675017, 
    -0.0546760970723012, 0.0149384047020821, -0.00891247040348825, 
    0.0102265252055527, -0.097934480213588, -0.0278339810388928, 
    -0.100665165599188, -0.0822709253417372, -0.0295680590569893, 
    0.00890200400941334, 0.0698881498430277, -0.136938054369718, 
    0.00102708191080007, -0.0183136686996089, 0.151645522891889, 
    0.603367255790234, -0.0679027553065585, 0.320500901701592, 
    0.587527758317801, 0.0890038543729782, 0.159648145356442, 
    -0.308844534434108, 0.107438958653252, 0.574480178287919, 
    0.304395749692516, -0.106292505145518, 0.43256983856424, 
    0.351678530391538, 0.118809373473583, 0.133652936004913, 
    0.352762118595948, 0.0341151454089076, 0.267146442009028, 
    0.687518529618163, 0.114333018874107, -0.0708820080320965, 
    -0.0282190909136195, -0.0329026947291645, -0.0357213283390608, 
    -0.0308990510265978, -0.0356930650685524, -0.025858579331519, 
    -0.0443363647378386, -0.0144390271952448, -0.103815925129504, 
    0.318977035630646, 0.231980956039951, -0.201487252137661, 
    0.265691855167804, 0.384574133120612, -0.0109104118608517, 
    0.0713802190629789, 0.211092312161803, -0.220654756323583, 
    0.642671939123754, 0.186382057901681, -0.0995406848621706, 
    0.435074743454693, 0.406333389220226, 0.211666265975063, 
    0.311803219128195, 1.14640756776127, 0.0553400486158265, 
    0.0739463003343155, -0.0222600514476174, 0.254877885184069, 
    0.352930258015849, 0.226181779663302, 0.164480844307134, 
    0.142119067227017, 0.118870325242182, 0.131389513777891, 
    0.129562219943938, 0.0560893609664141, 0.199445811085967, 
    0.292060192295574, 0.0959811620803942, 0.0833003707918411, 
    -0.202228096315254, 0.285774523488134, 0.254116650684332, 
    0.268115103369218, 0.580067950696886, 0.230525771442957, 
    0.111556313031154, 0.246511193626678, -0.149523981464401, 
    0.643028057444353, 0.429539609706873, -0.272543489043696, 
    0.272701673928159, 0.97770019660595, 0.360942124053235, 
    0.198265982738943, 0.765123620561211, 0.33367854676153, 
    0.0890084736395746, 0.0077853332265086, -0.0961299048711559, 
    -0.0746021946532451, 0.235533928829821, 0.0617502136901321, 
    -0.0683563365769856, 0.134123330174427, 0.0913464100333103, 
    -0.0455630201272065, 0.0109364066838505, -0.0561873710755185, 
    0.153822125467827, 0.0621864526591306, 0.0334588206320314, 
    -0.0390619517862307, -0.0405779889945126, 0.0780593646679777, 
    0.124979421792347, 0.0811624100750594, 0.0122801745013309, 
    0.0790758958517328, 0.129557759121492, 0.0734887581828975, 
    0.0460923781374912, 0.0994306079530748, 0.0896893969900539, 
    0.0646228173833323, 0.0448024780204084, -0.0789198755115377, 
    -0.0188370498752799, 0.0178271882362911, -0.0208357595194332, 
    0.0823757126719669, -0.00412566109616552, 0.0452364467397192, 
    -0.0170123301510371, 0.0309670426289482, -0.0551171126736989, 
    -0.0192967840185546, 0.152814579672137, 0.144304317939539, 
    0.00677891863434299, 0.172522136343696, 0.283371464020187, 
    0.166009588173607, 0.05100610965387, -0.0553181252452323, 
    -0.205548919687798, 0.353263051917109, 0.400213915592855, 
    0.266717697494167, 0.166424499502938, 0.118892434483146, 
    0.469837743065698, -0.205778865385029, 0.361541161062151, 
    0.860076094750211, 0.0548325960535258, -0.0813204062242369, 
    -0.0120096052833721, -0.0673214119615655, -0.114495347269221, 
    0.237560631660167, -0.0914859751076899, -0.0164492062961391, 
    -0.107957897018547, 0.1936803013563, -0.031480137707038, 
    -0.153353955705359, -0.0106933501867393, -0.0243825508435802, 
    0.00282219771344314, -0.341185553967214, 0.00101371885555475, 
    -0.261048481792244, -0.277004370095284, 0.170763524477354, 
    -0.323381221785649, -0.00721100999526154, 0.000485049100544158, 
    0.154967359455536, 0.168605009805453, 0.108782895122729, 
    0.0978452477663251, 0.0671612296310628, 0.144799051257436, 
    0.187301241231877, 0.114098214515914, 0.0976473919219449, 
    0.104690424074437, 0.0747968799262192, 0.10297351721217, 
    0.112584931430981, 0.120261817878252, 0.12634951339081, 
    0.165497486465994, 0.027634152383969, 0.0729262166261, -0.29596842100095, 
    0.550804720642022, 0.425250205849034, -0.097628573840242, 
    -0.108305106690304, -0.139405742266647, -0.261640948355043, 
    0.245688330362827, 0.70258421580751, 0.622349517179905, 
    0.134751264804852, -0.153449474151192, -0.122675863636596, 
    -0.0879626584906774, -0.00466377079884023, 0.0443530010715566, 
    0.0679525029449374, 0.0624905403354886, -0.100355409989385, 
    -0.0967215800159205, -0.229011871339089, 0.183938062726345, 
    -0.357570980807432, 0.0729297643649149, -0.580898569027513, 
    -0.167566372627391, -0.146826904060338, 0.0113294836552174, 
    0.216496218446188, -0.241193024859335,
  0.320592144948344, 0.748800023664597, 0.210633315061178, 
    -0.296610621988926, 0.292916616864104, 0.521350442054527, 
    0.136772350602829, -0.110609141648765, 0.307705760785361, 
    0.496505841916265, -0.330738626930482, -0.115602727052107, 
    -0.171330994170634, -0.0925376618600681, -0.113761523490396, 
    -0.0209580032044731, -0.23221664971539, -0.0470177703411221, 
    -0.228747143645213, -0.0780123879170475, -0.0982263349069673, 
    -0.0828848047757277, 0.0492009346473085, -0.0610227267319692, 
    0.121408908237025, -0.05801134568144, 0.0621897225333436, 
    -0.00865224590161084, 0.0630007013164954, -0.131029275606385, 
    0.00364646026290476, 0.0412587227259136, 0.0540470299578023, 
    0.0744478318647976, 0.0821236910047075, 0.0539845492722141, 
    0.0309899305783783, 0.0655716805979957, 0.159859746227432, 
    0.176120142329898, -0.0980430402719956, 0.256361455342788, 
    0.402971341952015, 0.169703249696254, 0.161457296908324, 
    0.311922820787626, 0.100805180931475, 0.145769569011617, 
    0.170546703005792, 0.445982872996576, 0.92787455070423, 
    0.543540554386695, 0.235184049703872, -0.421658236691624, 
    0.677802055103968, 0.842938807117005, 0.437278277411663, 
    -0.431436510132247, 0.48166808403227, 0.593882966054805, 
    0.0991509827365466, 0.0510024498143931, 0.406186785757626, 
    0.329311396298708, 0.106900479489735, -0.266107986839772, 
    0.154125087508393, 0.474086645700235, 0.0749260234999375, 
    0.0318432317243198, -0.202741015272875, -0.0666177120782027, 
    0.334571356068337, 0.426718453902199, 0.199832160044916, 
    -0.0608531833722682, 0.418343659402823, 0.20191895500931, 
    -0.172183319230534, -0.0203517236937459, 0.393657072329967, 
    0.303273531940568, 0.379780964529538, 0.183523444621541, 
    -0.0818846032292241, -0.203108357925169, 0.470195749058702, 
    0.133930339756399, -0.209037970481921, -0.0706580620644159, 
    -0.333029621079285, -0.0691914931683507, -0.038053364624738, 
    -0.20248180140175, 0.142904044277829, -0.164624826849864, 
    0.0520614824679094, -0.0807622992856322, 0.0378336148856223, 
    -0.218899571782732, -0.052463144073156, 0.137481520297496, 
    0.158709783324258, 0.0952796720241387, 0.263341033812559, 
    0.38035538840633, 0.207295791115463, 0.0573302783057729, 
    0.271145179144435, 0.420070811397321, 0.273574397219968, 
    0.182370748244887, 0.161323587620936, 0.176087052704241, 
    0.210562782965816, 0.187847235783468, 0.165591648735795, 
    0.193311978337687, 0.215001435238494, 0.187855872011473, 
    0.151543614828499, 0.134874772756916, 0.168509756777282, 
    0.224210876389356, 0.171642433803838, 0.0945170312444423, 
    0.22495573351813, 0.285546663047749, 0.141993705708317, 0.19273942078122, 
    0.321993386601313, 0.0869890186788082, 0.718135724141185, 
    0.421553669059204, 0.109841897343201, 0.0702957175330942, 
    -0.136839031695952, 0.0610068728119535, -0.200949577423876, 
    0.172725421985309, 0.88027495659615, 0.526937549926189, 
    -0.0189956548609205, -0.537781365918495, -0.104603717551393, 
    0.528919394416133, 0.242555559945175, 0.288897522136679, 
    0.487045129093196, -0.000451880062953408, -0.122108698311925, 
    0.0327548564498758, -0.501811983555588, -0.157701465737554, 
    -0.0324149622423886, -0.270147244558252, 0.0502834188531056, 
    -0.134659266443614, 0.027278917108843, -0.311903830486106, 
    -0.0554721984247375, 0.0501762518656529, 0.189304110345307, 
    0.32186158282354, 0.186203338676688, -0.15463736031023, 
    0.306653731512278, 0.559387393988844, -0.0225058598629176, 
    -0.152781269356476, -0.209808319365542, 0.510550617843696, 
    0.453235713641374, 0.145328181476685, -0.203757665010465, 
    0.0324713615177535, 0.555727257086429, 0.268499538715645, 
    0.0600400104646056, 0.123558527395542, 0.294574406949831, 
    0.31806454011809, 0.249979963525251, 0.196529720730818, 
    0.143131092537248, 0.158019277540995, 0.280880458562488, 
    0.218829652006947, 0.0796253184050711, -0.089038214615803, 
    0.345591376681801, 0.368598613529372, 0.0829045795676779, 
    -0.0589873508375988, -0.172210809277208, 0.368004703033478, 
    0.422550219234968, 0.104116023540321, -0.134080574410244, 
    0.0642964879075894, 0.393391555851374, 0.0529892040630738, 
    -0.0495564005628745, -0.139333223554403, 1.04876088779092, 
    0.0409450580009525, -0.412467796953228, 0.437754753996649, 
    0.401384536227915, -0.322407751123435, -0.179140201074861, 
    -0.0902737247281434, -0.147172117803067, -0.0213128985486965, 
    -0.173905125240898, 0.0226104449733013, -0.213552771831814, 
    0.00840667554894321, -0.193066442106673, 0.0215969517500621, 
    -0.137119824657894, -0.0153478270227744, 0.0606491963242488, 
    -0.0836548625558757, 0.0921443818347922, 0.0214261934990275, 
    0.0564434494790675, -0.0420078726620148, 0.0224596505354452, 
    -0.0892615983833944, -0.038517129550585, 0.0299906624588573, 
    0.0614657427380751, 0.0640907874412651, 0.0399921535742251, 
    -0.00428272665379671, 0.108684710483711, 0.216862679973529, 
    -0.0237089450214233, -0.223783227686109, -0.346739703074541, 
    0.117266679169916, 0.709474605101597, 0.34083623514745, 
    0.0467729178503962, 0.619843437562254, 0.174778889423786, 
    0.2592565003403, 1.33159762695118, 0.169717570129738, -0.113634841484873, 
    -0.0539885787714121, -0.0616696252488417, -0.101645192673756, 
    0.0544206432357151, -0.0726399636816385, -0.0549498239327306, 
    -0.0571948398708964, -0.16184232742522, -0.0804829731379125, 
    -0.083964949351163, -0.184784295102777, 0.118676491182799, 
    -0.154329622957641, -0.064752055618377, 0.0244174609506586, 
    0.0691903586358241, -0.021289718476132, 0.128654173756346, 
    -0.0994659543701057, 0.0598256744053496, -0.0428810298380239, 
    -0.00276922230655624, 0.0849819074470224, 0.0630811327057242, 
    0.104787228284471, -0.269886272282639, 0.177188846700856, 
    0.23946079381684, -0.233416188943714, 0.303693544264369, 
    0.422922095565004, -0.131613716828759, 0.900675697164954, 
    0.739411435207777, 0.679113314325528, 0.412811317553534, 
    -0.426810642623389, 0.187272003790927, 0.570682354467432, 
    0.0729942354772885, 0.119247224033438, 0.584750439832932, 
    0.228609991980961, -0.0414388239496697, 0.323157193572958, 
    0.335593249449832, 0.0733156363138145, 0.198577300001988, 
    0.453611308911452, 0.0288812999613823, -0.034412993960953, 
    -0.0620403856679582, -0.0626785267431438, 0.0403145884245014, 
    0.0435429816249738, 0.0274423632476496, -0.0140689721901469, 
    -0.0784156380378515, -0.0150395151169765, -0.141926777259532, 
    0.0190413016444415, 0.207254248998917, 0.413791990763701, 
    0.191266181704006, 0.00646494423847041, -0.161548539753434, 
    0.379739476667521, 0.261755376067997, 0.0388907373453198, 
    -0.0804638679641935, -0.0714921282788391, 0.0159768948736328, 
    -0.0843651086664683, 0.0124887730722826, -0.0634904327385104, 
    0.0104767759754036, -0.0157784686160963, 0.0746120277608027, 
    -0.0698838068357138, 0.0299223705417337, 0.0857845759639273, 
    0.109112456549361, 0.0954144127788249, 0.0904370651465937, 
    0.0909816657531822, 0.094858481374107, 0.0876733249771657, 
    0.0822772281006777, 0.0629069847849593, 0.112952245586184, 
    0.134492572612603, 0.13406427900078, 0.130234577862511, 
    0.140740341564144, 0.138577856017044, 0.12499991872304, 
    0.131408964710782, 0.143885812720669, 0.183976887428754, 
    0.185703657470829, -0.0255103557013633, 0.269067105959063, 
    0.339135114443045, 0.123820595650632, 0.163386881288462, 
    0.471719308542481, 0.483538924307383, 0.228810832170849, 
    -0.389048459771458,
  -0.0227653528852738, 0.0724890556245385, 0.1974960543363, 
    0.223445018453423, 0.128126652551801, 0.0247157660719251, 
    -0.131644096719789, 0.272829191410205, 0.429638371920084, 
    0.182855818710619, -0.12563036955727, -0.133491505343015, 
    0.874406766581192, 0.316683465484152, -0.324978746808187, 
    0.346029294513877, 0.618090759106283, 0.122564819727293, 
    -0.00240682281368071, -0.0118121859518007, 0.506361675901504, 
    0.0758928759647238, -0.0264466959182933, -0.0579485868776925, 
    0.147169958635781, 0.210545669691012, 0.11396968950593, 
    0.232729058512172, 0.211850148448323, -0.149347410484402, 
    -0.126172395212939, -0.166143589435941, -0.0364254707493362, 
    -0.285631290881585, -0.122796764240701, -0.131425872456622, 
    -0.211533561211652, 0.0577628224387352, -0.229638388055546, 
    0.0651990746705018, -0.126650446987309, 0.0440366421891637, 
    -0.0956519461326963, 0.0355159165604234, -0.0917590432588539, 
    0.0173208185916782, -0.125408663167758, -0.062181253424892, 
    0.0596973219423259, -0.135769219644621, 0.052953076601179, 
    0.0577400195586504, 0.0673103098658255, 0.0716896328194083, 
    0.0778678448961348, 0.0791525925737925, 0.0833241066336498, 
    0.0768282112118669, 0.0714613429881886, 0.0380310472919074, 
    0.0798972806798997, 0.118536894429636, 0.113335247527755, 
    0.119357834184373, 0.17225181494697, 0.133201982396871, 
    -0.0402209368926744, 0.29531625348267, 0.290408487801567, 
    -0.125716740198284, -0.0775401609291886, 0.429802517925479, 
    0.64726136154651, 0.289281680279307, 0.0207529747665718, 
    0.284514342232393, 0.0451529235440161, -0.043187921288721, 
    1.02675092612413, 0.411353465191983, 0.0199781073936803, 
    0.041061234588032, -0.120341608707425, 0.0172905002628166, 
    0.0932242780431108, -0.0074237754489236, -0.0297307345268055, 
    -0.0216833771436321, 0.232303704047237, -0.0815587957047152, 
    -0.214255539762699, -0.031680287236631, -0.330440461306788, 
    -0.107649022512858, 0.00910504897733065, -0.304274955554601, 
    0.0916450929971538, -0.0570470763739819, 0.0833595613136268, 
    -0.27821099385669, 0.104108816974552, -0.0205484938530157, 
    0.118749296255703, 0.321339659344472, 0.122675009005079, 
    -0.00707769420926373, -0.0999350453885034, 0.348629062675316, 
    0.316046400596175, 0.121493798509147, 0.0493709276292723, 
    0.0624416468572693, 0.453878448312783, 0.361483561444094, 
    0.0590540814371242, 0.109724520944738, 0.772787126959858, 
    0.504757934333518, 0.134861014099482, 0.0336444298109702, 
    0.610350007068421, 0.433212465196744, 0.109162209504102, 
    0.0983079328468584, 0.526188751179262, 0.259092608813247, 
    0.0417989066931248, 0.436418961703398, 0.318501400473532, 
    0.0289350159262624, 0.0284696059842041, 0.503621515336732, 
    0.254621366273521, -0.0391459728748609, 0.432558837953796, 
    0.411129593643519, -0.0854106986904263, -0.034783203236529, 
    0.0626593313739301, 0.517635123815977, -0.0434248503770975, 
    -0.0169341573345129, 0.0270602598677735, 0.145163125269508, 
    0.020926705875517, -0.0922636918021211, -0.12244860338427, 
    0.144244699036641, 0.194216810703353, -0.128804224964931, 
    -0.233237975203762, -0.0450582045426436, -0.287537136817343, 
    -0.185487070452579, 0.0898916105949446, -0.18455947085047, 
    0.0875791143102321, -0.127577793646618, 0.0450504768660778, 
    -0.262573349554167, -0.0169315499236562, 0.0387527122761708, 
    0.0761069339032538, 0.11000205963775, 0.121633750426824, 
    0.0898212686519335, 0.0922373269404806, 0.14620702765526, 
    0.115574213279046, 0.0470417422182276, 0.110203387041823, 
    0.17158638696969, 0.206831125785772, 0.194267938961681, 
    0.125994475591204, 0.0870253316408084, 0.346273541752562, 
    0.356280432537369, 0.0168309091948175, -0.102217033523108, 
    -0.251814131243336, 0.436118357814067, 0.395550493008011, 
    0.126910686579062, 0.0589177858846179, -0.205131405260857, 
    0.293020385947605, 0.167367007373131, 0.407134759239489, 
    0.785461113639943, 0.268201459859357, 0.103502216242574, 
    0.0926316138437933, 0.155820709543126, 0.436935535750167, 
    -0.232113923614226, 0.371967902022551, 0.65563332049034, 
    -0.0525105799405112, -0.0398933159977539, -0.073581336508228, 
    -0.243375855506376, 0.0412796652099934, -0.301218066848793, 
    -0.0391234979867128, -0.228343018932306, -0.0359644594974402, 
    -0.204178023821183, 0.0131850372763616, -0.215596672341442, 
    -0.00705363809755291, 0.0705974321186442, 0.0821633783354114, 
    0.088677586489105, 0.120863533449397, 0.101514999835331, 
    0.00196007232209876, 0.159819942748508, 0.139912589546204, 
    0.0494743834011679, -0.0927000900106398, 0.485731939489945, 
    0.194499300089254, 0.00745590551938377, -0.308846097484109, 
    0.326950841250498, 0.598646665875784, 0.118215622619084, 
    -0.041008683108763, -0.110852313487752, 0.223676845807622, 
    0.341554526174744, 0.143358075078609, 0.185792236074598, 
    0.311500148453905, -0.138053938982598, 0.303915369572923, 
    0.32025196295884, 0.102808885424811, 0.139076128219362, 
    -0.286487436465225, 0.0407796185428851, -0.598690598571217, 
    -0.231038666701474, -0.0522024698037759, -0.143025617295537, 
    0.0755368001253814, -0.300286114028395, -0.0311055510743786, 
    -0.347277644364948, -0.190512265140824, 0.086328291310051, 
    0.113907888951337, 0.100281557109047, 0.160020342307511, 
    0.175400578544439, 0.161069793660399, 0.170542050622332, 
    0.100757424506186, 0.0648586198739076, 0.120071323202969, 
    0.136207471627148, 0.162863705883, 0.20854393527794, 0.200600380100818, 
    0.137772182915989, 0.177587789308606, 0.33463585659907, 
    0.197974344588815, 0.00631676948539156, 0.174596177540248, 
    0.378410424289899, 0.050244762572846, 0.107567938237555, 
    0.627523557202394, 0.509363627173011, 0.328870054788996, 
    -0.0471703658855038, 0.629238320550415, 0.105580350200421, 
    -0.221602010005282, 0.139647525332691, 0.532603180136287, 
    -0.241474050020724, -0.616770353878401, 0.162488293935013, 
    0.372936329384961, -0.152878647095978, 0.0985495434280749, 
    0.0859157548599898, -0.134523640054696, -0.279548698082311, 
    0.122045043482721, -0.490621016490273, -0.07016492644094, 
    -0.365235964163595, -0.286475446624123, -0.175912943257686, 
    -0.258051062395053, -0.226472956616881, -0.0306883274456318, 
    0.0641279940814285, 0.156749870104664, 0.127269065272, 
    0.0598640682009727, 0.111361210018627, 0.00220456761747796, 
    0.0211675075147972, 0.112917040323663, 0.027857715369635, 
    0.199554442255823, 0.157888160934328, 0.0804648703729549, 
    -0.0200443608534263, 0.314600885543579, 0.223549165373835, 
    0.012896366810929, 0.480312030418466, 0.237449424279961, 
    -0.165108270508948, -0.152656817170713, 0.660482299475677, 
    0.354787275984668, -0.0294560660348271, 0.203185415683646, 
    0.931036141535932, 0.0474663101755423, -0.250126616818805, 
    0.473707922369098, 0.398191074656646, -0.299380036961928, 
    -0.12267562132384, -0.0315314285727962, 0.0723324663650405, 
    0.00950076692516208, -0.00852977317783213, -0.0670030589581097, 
    -0.0411923307292278, -0.192778317470399, -0.159700115839978, 
    -0.0224495969105222, -0.144722914422636, 0.0220339443100758, 
    -0.159462528081605, 0.0352362672566416, -0.158855344779064, 
    0.0185134773038846, -0.115938043202831, 0.0342640323001614, 
    -0.0985929221209591, 0.0568253872388326, -0.0333466618886109, 
    0.0106081430513401, -0.00530734567064531, 0.0168088946732381, 
    -0.0335592643797749, 0.00360111334802762, 0.0119546747444567, 
    0.01535234879119, -0.0546924623175452,
  0.275911518511929, 0.149059920282985, -0.032710754886362, 
    0.0966463547351561, 0.40408159841333, 0.228066575888076, 
    0.166559490243792, 0.475982317447487, 0.199771959710375, 
    -0.190722770612108, 0.0767495273490405, 0.57288540606839, 
    0.438579108951951, 0.211279079635595, 0.0666504109333358, 
    0.153805100074661, 0.14729875832903, 0.600709912251519, 
    0.403525021128515, 0.0456686759221393, -0.0474101934682606, 
    0.273602036154348, -0.213695371938986, 0.183534046990749, 
    -0.22813289152177, 0.0976810948958874, -0.214672862711939, 
    0.0507257410030891, -0.334598180913449, -0.137944664832243, 
    0.0154392857888215, 0.0261344864160265, 0.0348060530699078, 
    0.0948583547013391, 0.116215689080752, 0.0840960564196573, 
    -0.00359302204976469, 0.0456787119383904, 0.0657904317475004, 
    -0.00665302910640618, -0.0014486794058387, 0.0817654513233543, 
    0.098904500975281, 0.0654120502199129, 0.0394659958772666, 
    0.105069728920371, 0.161045654269688, 0.0779488579076004, 
    0.00215199502574756, -0.2112252411984, 0.12235599844154, 
    0.721340439033924, 0.217900841531642, -0.215889183302904, 
    -0.298738959895602, 0.409903656239259, 0.644532887248805, 
    0.173471527396049, 0.0246228584604686, -0.216324897987236, 
    0.231483428460644, 0.235918138756991, 0.210916755501681, 
    0.643336600397772, 0.227170620438281, -0.33614967197305, 
    0.399588321109843, 0.320570348357964, -0.0496397499856914, 
    0.129673182422494, -0.468354678319698, -0.0288915320476687, 
    -0.232459267535602, -0.308114520858801, 0.146184114287682, 
    -0.310469954591504, 0.00365394555742535, -0.1001494536749, 
    0.0180188707138642, -0.328611522141601, -0.116939646233252, 
    0.174952346731957, 0.143182103592185, 0.0779596236014538, 
    0.0530562035818629, 0.131291347788207, 0.0430489361972514, 
    0.233925429757819, 0.522791189542633, 0.103689542044973, 
    -0.137164175760632, 0.139214192707445, 0.566115840061826, 
    -0.0468472657894532, -0.259971771299626, -0.156576944494412, 
    0.646297690449782, 0.417070852675054, 0.347036571480255, 
    0.552923909178537, 0.126708215780783, -0.0170296543110631, 
    -0.0335029435764813, -0.0613871167832895, 0.00526878205447147, 
    -0.0437785488662644, -0.06014472785214, -0.0241704620969012, 
    -0.0514652601303396, -0.066784172804172, -0.0730376151046492, 
    0.0332194731923513, -0.0325346769138407, 0.0278910723924226, 
    -0.117764548451133, -0.0160946146408995, 0.00236207128982591, 
    -0.0265461867968512, 0.118391635954242, -0.0796482137228157, 
    0.0519816920283742, 0.10652461865966, 0.0412363299748969, 
    0.174956166235243, 0.182173946427347, 0.0270931975824429, 
    0.142892227472481, 0.309976958832261, 0.0925463576913717, 
    -0.110046031940453, 0.236454554672796, 0.216485499787655, 
    0.395072819904507, 0.654889563864566, 0.101730113096401, 
    -0.02234575570914, 0.284764357690981, -0.591309290539322, 
    0.625005745457468, 0.701683401776781, 0.0270615099824711, 
    -0.0400314308789605, -0.269112086277424, 0.0377811172923287, 
    -0.0483375040149741, 0.621903682711108, 0.00225377623915308, 
    -0.0975326291302371, -0.0652440079309417, 0.0229380400414326, 
    -0.469101707994495, -0.218152805232032, -0.00912831810266142, 
    -0.262328518453387, 0.148895093669576, -0.213326752735647, 
    0.119730736640817, -0.138089836789861, 0.0940786907605334, 
    -0.311230448398623, -0.0287414126120099, 0.0862113838099988, 
    0.0643969220256471, 0.147442232229083, 0.244063719441795, 
    0.124205851858843, 0.0621496267352026, 0.330776953784844, 
    0.42808198684697, 0.270388166569905, -0.258896296874789, 
    0.622504270909763, 0.373467219573116, -0.123806503220785, 
    0.22404332297074, 0.768182843930325, 0.144051961578474, 
    -0.347780795666207, 0.305617011210356, 0.643464512369907, 
    0.121928227792471, 0.000632939391219584, -0.00897758483369013, 
    -0.209400262604158, -0.00863789777040065, 0.0174826173557642, 
    0.424015848712318, 0.439788686044717, 0.386014083086669, 
    0.323096853202843, -0.110445210630981, -0.227557172856729, 
    -0.136153556639422, -0.154457690139392, -0.136917588596863, 
    -0.132279898311209, -0.113980643165777, -0.0708116448705374, 
    -0.166939239796437, -0.190791010355873, 0.0576478661204361, 
    -0.0440877337877211, 0.0390123040082309, -0.0362012580340706, 
    0.000940609078301125, -0.0449613077223911, -0.0728112252295545, 
    0.0429155742483102, 0.0522010422959837, -0.0514604926292117, 
    0.145490856125323, -0.0865047910248999, 0.08107272037577, 
    0.460860635947127, 0.0569037555287973, -0.00587025240933059, 
    -0.0446460994338454, 0.412641983480746, 0.0704086656087668, 
    -0.0244889739835412, 0.0758214101369431, -0.117676184030945, 
    0.0106297500769684, 0.920675086668945, 0.197475706862307, 
    -0.109644390042074, 0.0384606198834341, -0.275114525694458, 
    0.642185232571526, 0.0873169526770174, -0.110633674420389, 
    0.0749154253517679, -0.0783066627199809, -0.00143782813461749, 
    -0.334361071775989, -0.0813181254106939, -0.0441152822082559, 
    -0.0412612289872257, 0.119635319558552, -0.239053761893676, 
    -0.0170347911841525, 0.128790422291892, 0.124391705949564, 
    0.143017168083291, 0.2404718026845, 0.251477890469619, 0.252384514109508, 
    0.274729503293424, 0.181029436621649, 0.11595062012084, 
    0.445181386928745, 0.37811480594317, 0.108201001248029, 
    0.0815395648635502, 0.586778987037675, 0.308517849902446, 
    0.0418736942382061, 0.59711777322625, 0.383257686151562, 
    -0.0262863696583623, 0.389514582931954, 0.576795651452512, 
    0.0514130325376394, -0.072179498988956, -0.162419781902313, 
    0.260520148117019, 0.552171048031074, 0.313867309388471, 
    0.0701195461173609, 0.0757440767746052, 0.623320231262235, 
    0.208548191396899, 0.039465470824702, 0.0347528878747871, 
    0.0501214871074722, 0.202267418369117, 0.0593220201809009, 
    0.522891566459525, 0.185839614407718, -0.0582480866467603, 
    -0.11443063260053, 0.0318828638443722, -0.115056035322234, 
    0.0147605604035274, -0.234222549573284, -0.0593481469002818, 
    -0.0607839519480458, -0.131989079776755, 0.0899134161717389, 
    -0.168116847824705, 0.0834127428619694, 0.0520963184807725, 
    -0.00145442239572556, 0.350163163495177, 0.240799240620822, 
    0.0506578251364456, -0.169044578215291, 0.175629861939618, 
    0.489428947920135, 0.306471958830687, 0.120602033322822, 
    0.735099600995538, 0.180284017052406, -0.0609301851436124, 
    0.0841791577910652, 0.873684568253744, -0.0986563911781064, 
    0.00430943803926831, -0.192735559501872, 0.663173919357142, 
    0.257319400806503, 0.100102766120245, 0.0574203504018468, 
    0.231883122854177, -0.216424256680661, 0.519007905655205, 
    0.433821408404907, 0.0552913014492207, 0.33484747554674, 
    0.535993398278969, 0.197238699737455, 0.0945273310848065, 
    -0.0654033316698912, 0.222343015543172, 0.0691632847825943, 
    0.0452294106982636, 0.100147623093277, 0.00175460418281842, 
    0.181889018469484, -0.150843765087177, -0.171573160486348, 
    -0.107538992933443, -0.0767920249203021, -0.119491310197548, 
    -0.0643857751082946, -0.0848861123774335, 0.0224524119100761, 
    -0.131759207484126, 0.0786264790685549, -0.107833506453537, 
    0.0442091729059651, 0.0262121538957002, 0.0664443712412994, 
    0.00866516992766243, 0.063959863822203, -0.0253915536306586, 
    0.0308460462374165, 0.0216280425959885, 0.0575809998819131, 
    -0.037920227389759, 0.0367043740804994, 0.0734721512418959, 
    0.0905404507712644, 0.0968170372509932, 0.0971327459989401, 
    0.0891536279020188, 0.0973739230728642, 0.0917037533871209, 
    0.0497245075147737, 0.0592716184672001,
  -0.0280583583481647, -0.007706193629905, -0.153583670935259, 
    -0.0189787800685309, -0.150385909478643, -0.115136188547608, 
    -0.0197980665455689, -0.0427477221395905, 0.0101075155830566, 
    -0.123058811523574, -0.0250026065350413, 0.114412777298092, 
    0.235561743424868, 0.174831268611454, 0.0967493769069186, 
    0.209139252261334, 0.408553259957002, 0.330819069449916, 
    0.156003693759204, 0.166426319573121, 0.505566933699488, 
    0.324750925906981, -0.00635196411981887, 0.383953825058978, 
    0.715160967274405, 0.244891391906292, -0.086449841363114, 
    0.427069410499818, 0.553493191554388, 0.297395567130541, 
    0.153568142322857, -0.0607080517257681, 0.16453877752083, 
    0.603361669250226, 0.212144359030998, -0.0332205204292783, 
    0.779819530798443, 0.570341888602756, 0.19317863385501, 
    0.0355917451208349, 0.170825274630773, 0.42874038706901, 
    0.127119264126774, 0.214742621908921, 0.12811024180333, 
    -0.225142501214946, -0.0581824229873773, -0.0352669726203133, 
    0.110705545444867, 0.371753647803868, -0.0823833714577017, 
    0.0048133002563084, -0.182417638729592, -0.0172917525660078, 
    -0.154931583894083, -0.132283143141565, 0.00358832401191836, 
    -0.0795909450968982, 0.0644597133330903, -0.161767558402628, 
    0.102051651589293, 0.108690169835763, -0.00192034229717833, 
    0.447867272943815, 0.223678066933515, -0.0025681363852894, 
    0.0557702532830274, -0.247898819613862, 0.719147188652233, 
    0.295631125626508, -0.0667694778182779, 0.321842699357059, 
    0.407825039914409, -0.047310216185279, 0.58472884482641, 
    0.899430298811632, 0.453182542056613, 0.0949414037457065, 
    -0.123023140764382, -0.0963085864193067, 0.595707283010701, 
    -0.0757320907309335, -0.132285855290137, 0.125587786026849, 
    0.20646066300489, -0.173231565795903, 0.0151542880697304, 
    0.461645913593366, 0.195038994722064, 0.00471135380219449, 
    -0.161746467809504, -0.0402661916546636, -0.159572251223293, 
    -0.151779058241249, -0.204584229239265, -0.013435381087493, 
    -0.188630771626016, 0.0603266482532581, -0.179824135987627, 
    0.0597981169747614, -0.107993955951131, 0.0141181490725214, 
    -0.109382510993807, -0.0194697513228559, -0.147562943054451, 
    -0.108651623633629, 0.080054939640343, -0.0593667928803069, 
    0.152723411051882, -0.0793809968089713, 0.368316883945158, 
    0.166849859781348, 0.0278040002318092, -0.0448498373355011, 
    -0.0999919937149778, 0.349235279819954, 0.508737667682359, 
    0.0462763051977614, -0.176914089822886, 0.0227330982765003, 
    0.536260058297332, -0.108984801461677, -0.0208099826482005, 
    -0.429165327810489, 0.521227180391138, 0.532657445655295, 
    0.185500496091665, -0.23584741856014, 0.148213672138995, 
    0.454283265915312, 0.217733808876151, 0.325270973018293, 
    0.322360463074935, 0.104469181228614, -0.201847153896444, 
    0.411028882437354, 0.445831470758146, 0.0741064229550383, 
    0.0179715745434487, -0.131326515822052, 0.310823526666076, 
    0.242105333399448, 0.278403929022852, 0.209058774984974, 
    -0.181193424426125, 0.0207235002203531, 0.50839836361101, 
    0.17501838064754, 0.0706392317308716, -0.0253767903719408, 
    9.41185742336787e-05, 0.175710912707296, 0.111537237398211, 
    0.139537737900628, 0.367829128051282, 0.360874327044099, 
    0.27932627144791, 0.171777204954128, 0.0401404271856816, 
    0.079421173046378, -0.174972393997642, 0.13777940789849, 
    -0.242991039339399, 0.0512922113132687, -0.270776627948799, 
    -0.072311426643369, -0.270259644935462, -0.180720470880079, 
    0.13054933500087, -0.324394073202047, -0.00453060187266578, 
    0.0838159197816806, 0.0761825897555532, 0.123675419227435, 
    0.1513565335084, 0.111792331605336, 0.108260119818713, 0.176026188512807, 
    0.135253118132129, 0.0171368890302009, 0.189854328732609, 
    0.309784758713128, 0.145842870107834, 0.0361192760849402, 
    0.482734653222812, 0.319073025625411, 0.0654118192366384, 
    -0.0219622905080517, 0.457635861923153, 0.405110721571675, 
    0.248242245908205, -0.237663328925291, 0.365216437212558, 
    0.482746111058314, 0.126611151173234, 0.0354076230396275, 
    -0.310645744715617, 0.192800167124775, 0.615232214409522, 
    0.0657981228724874, -0.125507512743721, -0.0979031909957761, 
    0.361370586618211, 0.145930577049043, -0.0518748561443559, 
    0.199964066973539, 0.406455243204144, -0.0421639412960999, 
    0.34910894248624, 0.380420808060519, -0.183946140235217, 
    -0.0649189748355462, -0.11154191163829, -0.068343809506616, 
    -0.0294556429447095, -0.0682754228463122, 0.0508860423513154, 
    -0.0359236673275806, -0.0475494365893641, -0.0201140872254749, 
    -0.0252119797745316, 0.093614701765544, -0.00321477998137797, 
    0.0836044249077387, -0.00437773451201887, 0.0811068822126179, 
    -0.138584415843396, 0.0352564072777664, -0.175351530961194, 
    -0.0766068767798234, -0.0163322315117091, 0.0546442037328381, 
    0.065067206293937, 0.0717869092800119, 0.0694320526223475, 
    0.0694013208891677, 0.0535198125108396, 0.0601020156966879, 
    0.0435647143907855, -0.0124011882474813, 0.0877619824616639, 
    0.122552997950725, 0.144086091911641, 0.181075815032683, 
    0.22884085150494, 0.248714499751655, 0.132281791774955, 
    0.0653056016733038, 0.500560055717429, 0.188392384462875, 
    -0.00959242368782448, 0.118379930281567, 0.59214159714756, 
    0.0942953760261424, 0.139097535897896, -0.275362107949054, 
    0.559274118247957, 0.297586533896481, 0.0767920576393398, 
    0.262728480537624, 0.235520876576712, 0.0402697867513233, 
    0.0511271364736774, 0.103100203783859, -0.110090644396132, 
    -0.0406336656629917, -0.0795743610274002, 0.0719786103474896, 
    0.0044233229095941, 0.197314852796106, -0.180017051955548, 
    0.184857246640279, -0.16964040772938, 0.0975449765254842, 
    -0.0318506469277166, 0.192260135013981, -0.249989927282774, 
    0.0933308624521856, -0.467537262400844, -0.178839879523713, 
    -0.0444897145290339, 0.0272951032789341, 0.0944066130433278, 
    0.115239811007301, 0.111231905219192, 0.0686632751505178, 
    0.0624734821980442, 0.167704766983267, 0.156786202369881, 
    0.143557360651184, 0.209890669553502, 0.0359145144557579, 
    0.149472386688785, 0.572189276577901, 0.218957358147274, 
    -0.0378799616285803, 0.014672785600199, 0.490666755259699, 
    0.274070484984485, 0.374644990190732, 0.374663721122925, 
    -0.214037312210438, 0.307085467177519, 0.520170078424296, 
    0.143867166062461, 0.163767780090392, 0.166329424658807, 
    -0.190464176685309, -0.0798414489020566, 0.704323034892833, 
    -0.00986857485038223, -0.0518065271493571, 0.167733740544224, 
    -0.120735016590579, -0.281421671852224, -0.0347247582547649, 
    -0.0993466300584494, 0.261359385127752, -0.0939210300418268, 
    -0.0881221984802472, -0.244709325364709, -0.190251722333271, 
    0.0518638767499933, -0.190010138924289, 0.0993753355325582, 
    -0.148818676661952, 0.0838862082888466, -0.0973389379430913, 
    0.088132347860219, -0.217525743987298, -0.00185692564452235, 
    0.0621269834772026, 0.0915364562880648, 0.10882637794426, 
    0.11498636457179, 0.0824748471085812, 0.0755916764733234, 
    0.159973599646001, 0.12075967786705, 0.0339405504306766, 
    0.0740622649642635, -0.111262425274511, 0.392840925566096, 
    0.360585826617331, 0.135056927506925, 0.0269070769075737, 
    0.319054947906228, 0.353030178825081, 0.0668560542590643, 
    0.117943269170756, 0.863835746912239, 0.0823262844045438, 
    -0.0408210685350421, 0.240928214849796, -0.309203447652957, 
    0.302440436710539, 0.178427223262405, 0.0928665884899219, 
    0.902322387749399, 0.338101542208183,
  0.0989637053959037, 0.0105598492439582, -0.158807298654518, 
    -0.124466393324318, -0.118672867782682, -0.113560317738941, 
    -0.189496315946423, -0.163534269817934, -0.150749611129717, 
    -0.0769362593585187, -0.162891656546721, 0.0705564793519466, 
    0.285160790396987, 0.162053758229591, 0.0623037307456755, 
    -0.0655842366061423, 0.180682270274123, 0.435036802620751, 
    0.134611111152205, -0.0310871012243959, -0.115006865009383, 
    0.212303350982943, 0.481918163310003, 0.213181529912466, 
    0.165120116445283, 0.318278918658464, -0.172171868545746, 
    0.252163938823562, 0.51116604815609, -0.0670024350958659, 
    -0.148445306553357, 0.0322388635851206, -0.167942503408738, 
    0.0283705591981164, -0.158835493166758, 0.000859303609734394, 
    -0.252374927140784, -0.0594109294102259, -0.184058239499517, 
    -0.127890726433279, -0.0595348062712115, 0.109181274429799, 
    0.177390487290341, 0.148243411698875, 0.116088553534954, 
    0.143069748091718, 0.22950655310217, 0.220550771395104, 
    0.159214247769187, 0.146818489730698, 0.167555933242454, 
    0.176450190340359, 0.167884220598728, 0.140796119155872, 
    0.164733269759164, 0.246898618831542, 0.167556368383609, 
    0.014532421730276, 0.267866891028858, 0.249227357560433, 
    0.00146780902295172, 0.0649589400584573, 0.600933062649647, 
    0.319974547496121, 0.247527412584592, -0.229832185212361, 
    0.442613431237763, 0.389910053430106, 0.200249666816407, 
    0.198854497822755, -0.422514259737283, 0.441186327459082, 
    0.72760509416093, -0.2331411412354, -0.0338484683882289, 
    -0.535632491239709, 0.96011622921356, 0.262951609177558, 
    0.0105762140791754, 0.0119970761220351, 0.469644897092445, 
    0.354731648967677, 0.0957841578814539, 0.0112420888143857, 
    -0.0551497421132233, 0.281686478812178, 0.160411591978777, 
    -0.00548930506953688, 0.288385825540735, 0.20737255927137, 
    -0.065511342863515, 0.168146507544089, 0.485547830782714, 
    0.17272937182891, 0.0423985064489035, -0.0134338987726609, 
    -0.23240703944667, 0.553751482207339, 0.153342567537667, 
    0.0475860100942933, -0.163021867444201, -0.0350493458100217, 
    0.485322939444021, 0.256822042376706, 0.139511912201115, 
    0.175139669364999, -0.090174265449384, 0.274087248762587, 
    0.699203276069085, -0.146841501090131, -0.166363029556475, 
    -0.0952757291974416, -0.0548071952359149, 0.0174380511891672, 
    -0.110054397189648, -0.103043117080839, -0.0172909793534936, 
    -0.116970545180152, 0.0140131020410317, -0.100682542923141, 
    0.0663067713102917, 0.0644017633550853, 0.145219379414039, 
    0.207386261589265, 0.181192169165999, 0.1292773102272, 
    0.0837498798271864, 0.125040735677167, 0.226516775140445, 
    0.192853377540597, 0.0805325306452049, 0.0521208277746951, 
    0.0743919467274619, 0.0907152492388996, 0.0977204404052807, 
    0.0728568485447673, 0.0842449145781549, 0.0790644405905117, 
    0.0863723637666239, 0.0563374352313308, 0.0947388875277499, 
    0.107828710415106, 0.110960636480893, 0.111516413048388, 
    0.112353557242648, 0.0999061958751962, 0.0897069945100397, 
    0.136152801421186, 0.169215520214212, 0.0904021756418188, 
    -0.0220213001728244, 0.0568760990802525, 0.406678989398406, 
    0.212175902210219, 0.0215641707365187, 0.271114487846226, 
    0.284337230164779, 0.103500621430828, 0.608101381979201, 
    0.354111929556309, -0.0958691032095515, -0.221579936977999, 
    0.597698070831495, 0.833201574957013, 0.023670335322966, 
    -0.579060739707817, -0.0405686848862009, 0.99812096011908, 
    -0.086091435920554, 0.00180094483149618, -0.261645259228836, 
    -0.166503311389705, -0.184486319724928, -0.219427828693252, 
    -0.173760980855747, -0.0180697041488527, -0.11474414762769, 
    -0.353327195448876, -0.0333674993018962, -0.215983078563547, 
    0.027858163542285, -0.202448304100956, -0.207649999925316, 
    0.121412010751423, -0.0471089743020712, -0.259490534721806, 
    -0.00725430679109139, 0.0143656130955697, 0.021701249927708, 
    -0.321303990381493, 0.00146271622119484, -0.0802858980757817, 
    -0.04524336567084, -0.0784517859094197, -0.00866492332936475, 
    0.00324065774393306, -0.0613021668803574, 0.113130940194355, 
    -0.0224628075242173, -0.00763891282277157, 0.305030703375686, 
    -0.033130252316684, -0.458790738837959, -0.0776327777224556, 
    0.550614953210111, 0.443426058156963, 0.348431859862848, 
    -0.260315958135093, 0.912026207303981, 0.456863393900987, 
    0.0302065364358778, 0.0589922876918309, -0.0425944995397602, 
    -0.0168428150975626, 0.157940095731298, 0.088279253863667, 
    0.0789724872045069, 0.130883368699516, 0.223925040026014, 
    0.0736218850703422, -0.0169437231348482, 0.0229529250758787, 
    -0.0529823944189069, 0.0157656914539772, -0.0834781817127852, 
    -0.0281920336918705, -0.0265177386354751, -0.0343453780409161, 
    -0.0559381585406414, 0.065714050390252, 0.274263161294219, 
    0.00318106370579647, -0.185581125046048, 0.402144411503808, 
    0.355585851472431, 0.321585021445754, 0.275735937639303, 
    -0.208075506652017, 0.393089208503199, 0.378768784823591, 
    0.0957169388111191, 0.278493369885509, 0.360547915972331, 
    0.0604255627409877, 0.250397205903425, 0.468805127526214, 
    0.0961184257148289, 0.33537250974684, 0.692581358100615, 
    0.123515194651771, -0.0535974498531285, -0.0214761607661604, 
    -0.0144597368120869, -0.0231368628031232, -0.0194183780602782, 
    -0.00117479651596218, -0.050491082047836, 0.0410357607827205, 
    0.0377775464927872, -0.0726105262943414, 0.156613552599915, 
    -0.0702658252229833, 0.407361549643267, 0.298932267487098, 
    0.0873871300285677, -0.0884240931465638, 0.0836852829992371, 
    0.0352041361161861, 0.633196990243246, 0.391349467778948, 
    0.00339249357749999, -0.184348889696786, -0.20506470708709, 
    0.960038390272952, 0.188076594252203, 0.0893837383106746, 
    -0.250468672309631, 0.287955270257988, 0.435869088822493, 
    0.451935986757559, 0.532043227859058, 0.320993010794473, 
    0.115930100961608, 0.0679320696409951, -0.130508772999361, 
    0.00197492054438342, 0.234135891626424, 0.142729753930278, 
    0.0420448040046472, -0.0194413582112011, -0.0946919507813341, 
    0.253647415464192, 0.239613739115853, 0.115946683295779, 
    0.0746575770004936, 0.0793054482055444, -0.000600885336852888, 
    0.0925647158689075, 0.456766580631101, 0.230032248393528, 
    -0.160477529129853, 0.41931602711724, 0.474217817801917, 
    0.0749391209520838, 0.179799504074241, -0.121660373761005, 
    0.477394347325685, 0.238005505737254, -0.00488385242023953, 
    0.382213994707003, 0.234249365581003, 0.0588152893666693, 
    0.0115865866008346, -0.0160798846433334, -0.0210183815987301, 
    0.0106471568365769, 0.0168208227799002, -0.0498630405441006, 
    -0.0460411614200544, -0.0397024184573633, 0.0213103636348703, 
    0.0147572586920504, 0.0229284321707684, 0.0171826774233916, 
    0.0289406181862758, 0.0169488873859194, 0.0378570925686511, 
    0.0399762442219033, 0.0665125373463501, -0.00849098500882148, 
    0.0341721738860673, 0.135297905993343, 0.216031876832486, 
    0.149775779121661, 0.0429721267260714, 0.0519075428257893, 
    0.241111660862514, 0.433741011989588, 0.247628969598849, 
    -0.256419915898637, 0.26080705302811, 0.72679330588387, 
    0.256256998822163, -0.313616917733369, 0.28220953730756, 
    0.444230198888443, 0.155694579895166, 0.868320082467213, 
    0.477132243994276, 0.0249762324942048, -0.184089215248071, 
    0.750356758559441, 0.254875187925943, -0.00271895779376753, 
    -0.0658388278626228, -0.41164830667192, -0.319170630280958, 
    0.502105873343289, 0.484579553156257, 0.267500468221585,
  -0.0979601252361409, -0.114098897298055, 0.0925945446586936, 
    0.112302832396513, 0.0550751849064707, 0.0922591741658795, 
    0.258754169117347, -0.18873023705575, -0.182267861447322, 
    -0.0354057856169636, -0.228717748810721, -0.0855238522160879, 
    -0.208427361170087, -0.107575290673586, -0.182141284395541, 
    -0.144745968794662, -0.0861231358800177, -0.168336302119857, 
    -0.00469391864054092, -0.168585206638341, -0.0139196150056548, 
    0.0693974055311661, 0.0744483676359074, 0.0850049197851641, 
    0.0779325589283908, 0.0762744877900675, 0.0825298232354136, 
    0.120035223332357, 0.0812817742241581, -0.0689870598949546, 
    0.125275462522774, 0.261446076697689, 0.0705746710294032, 
    0.191118156836034, 0.461698919657441, 0.0873713859845505, 
    0.00594376307811954, 0.0357968149936071, 0.261121455157923, 
    0.0680391485372631, 0.557070841588459, 0.300170556953488, 
    -0.199990231448084, 0.0344283700816275, -0.348722648981882, 
    0.459517240494959, 0.11762504661027, 0.361736541191632, 
    0.985101279996245, 0.240224856497815, -0.0401897149464915, 
    -0.0268300613461796, 0.0597422454422659, 0.014637740023327, 
    0.0603951542109587, -0.0591456783842481, 0.0333065905360426, 
    -0.029055814444134, 0.0406889635395401, -0.061365966221688, 
    0.0826245497394697, 0.122752461650376, 0.0812128200767935, 
    0.113588495363993, 0.236673896574462, 0.260632361023977, 
    0.238187086525474, 0.194859491769507, 0.103692057793986, 
    0.245020789889634, 0.423298024640631, 0.166810971233876, 
    0.100389105384701, 0.742532378734688, 0.223514526821381, 
    -0.237948703293831, 0.192032616619286, 0.758714668877505, 
    -0.032885561618333, -0.0614217883958618, -0.300940716204413, 
    0.364346581283228, 0.617606632353405, -0.123077060673485, 
    -0.195745726429328, -0.358579030586366, 0.320447869390377, 
    0.48015106563641, 0.264446336564072, -0.0262989290839243, 
    0.287478473078206, 0.151789342825257, 0.002928652560741, 
    0.0475360079430187, 0.0708317527559727, 0.200846344494615, 
    0.142814215598828, -0.336536841469816, -0.408033358460725, 
    0.0159541234979689, -0.270009094105002, -0.136394591924954, 
    -0.0329232514937089, -0.204578054855568, 0.127676116494104, 
    -0.194889889333476, 0.0999210354007874, -0.216118395305181, 
    0.0410538389032142, -0.216703411186337, -0.029544346183219, 
    0.0643148853119095, 0.00577389663578755, 0.205649918872575, 
    0.195947182688958, 0.043866342353208, 0.029486483552501, 
    0.333586735538136, 0.0584900239149167, -0.00276128644775944, 
    0.368233501710162, -0.243960427153735, 0.777387080071338, 
    0.520827056437869, 0.055707527665649, -0.299240638843694, 
    0.0247480401619559, 0.658476016473529, 0.384214576283236, 
    0.145391039083701, 0.0886240127714238, 0.339003250279298, 
    0.130337665064065, 0.0899685943456481, 0.338056049115947, 
    0.113742112875065, 0.00241103494324819, 0.181504175633187, 
    0.119817717956098, -0.0366422532116323, -0.0738797540987357, 
    -0.0192645529502479, -0.0816111275766686, -0.0433299981620392, 
    -0.04444110079509, -0.0406634635365464, -0.0632638314280201, 
    0.0303665700797098, 0.0353361659522776, -0.105284861845582, 
    0.0224259665006119, 0.0204009347223736, 0.0572208731343564, 
    0.48717881801119, 0.220352729038269, -0.0894596426643802, 
    0.328349336539993, 0.318282817713326, -0.0582651218526887, 
    0.0627310257953707, 0.550898191999783, 0.0267140113890805, 
    0.49385645546708, 0.876643288338384, 0.537922731081668, 
    0.304365965506667, -0.199991805855925, 0.249021667171683, 
    1.18271428091656, 0.0945493037629938, -0.132666296127302, 
    0.0177735969374542, -0.184418071232912, -0.0655536562324167, 
    -0.0773558223132426, -0.117217369127656, -0.0739243224743784, 
    -0.089600059277715, -0.00653919065855699, -0.119051431336058, 
    0.0376414867735339, 0.0921447082492156, 0.102418240924344, 
    0.0920492488304135, 0.116746088615789, 0.135328529919987, 
    0.0835031958010405, 0.0231670151234982, 0.176572642395878, 
    0.221172048817021, 0.160207052024867, -0.167935720165937, 
    0.0117853958902594, 0.493324566986944, 0.528969654857368, 
    0.329617181934198, -0.267511123315322, 0.610181447751556, 
    0.386927563443975, 0.124526686766212, 0.727644075303734, 
    0.40893056481647, -0.301601102693448, 0.338110314398002, 
    0.548205343595619, 0.0936768469898271, 0.11618303484144, 
    0.114853219810919, -0.293681966887662, 0.440328376756098, 
    0.296564595435822, 0.00923131765566063, -0.0640723906433019, 
    -0.00726852667021828, -0.117641163994837, -0.00154023642473498, 
    -0.00064205156492235, -0.0187755358053153, -0.00914015201383592, 
    0.0241164942687738, 0.209746291143044, 0.0467787105287867, 
    -0.0472118735981027, 0.250138031249907, 0.406920321000038, 
    0.183687307698296, 0.0472153106873821, 0.077394424415854, 
    0.118583999994678, 0.136356146272896, 0.364320851542991, 0.3339901175958, 
    0.127644125101433, 0.00883480258445338, 0.237531225567875, 
    0.296598366336594, 0.139401403615254, 0.0897148393476024, 
    0.304791609966734, 0.200537208003082, 0.0309649443826191, 
    0.0152092652913436, 0.0511027130150678, 0.0503247612027486, 
    0.0616477974138815, 0.0282555847629529, 0.0380461486597255, 
    0.0886969342656046, 0.0720321697428286, -0.0254043238016262, 
    -0.0511542792924962, 0.258444667363253, 0.251810784673426, 
    0.109423089311055, -0.1371567226086, 0.172248800600506, 
    0.369449384892655, 0.133354549141996, 0.0483988256606222, 
    0.0274338464269519, 0.400870403863765, 0.068943537502468, 
    0.845273196476068, 0.441641724163441, -0.0537645664670706, 
    0.094926248754562, 0.676637672080521, 0.283230907104422, 
    0.362338485813436, 0.340184485518058, -0.214445322537634, 
    -0.128439698897158, -0.155283160502788, -0.115371732533524, 
    -0.194289539984707, -0.0903902218571571, -0.207236356017578, 
    -0.111385408189659, -0.175426901045724, -0.125542902011065, 
    -0.0675910823889802, -0.0394966030572673, 0.00685707961556083, 
    -0.085635451438861, 0.0853031897108774, -0.0127532585661488, 
    0.0484503894880785, 0.0104899650099094, 0.0497973926536777, 
    -0.102724584074938, 0.0331957851961033, 0.0873268498972096, 
    0.0582218291520921, 0.10899223289197, 0.180013003829972, 
    0.144006407520466, 0.14115283328357, 0.168306474890407, 
    0.0693436046159908, 0.0176183499960842, 0.493563920678272, 
    0.27744228801275, 0.0489541827261013, 0.201682863673367, 
    0.16921684562966, 0.142987727481944, 0.797165990755518, 
    0.431967207737629, 0.076349659161082, 0.655788029264247, 
    0.482189106728669, 0.351956129854055, 0.339288180307868, 
    -0.248307218640367, 0.212493659746977, 0.447353763615929, 
    0.370466578538112, 0.194111281534547, -0.00214402160130295, 
    0.00983013107414248, 0.379657515420704, 0.0618007641220154, 
    -0.0414583214494841, 0.201339688685319, -0.0153799958123559, 
    -0.123805822213155, -0.152315405794507, -0.0869873622013735, 
    0.0875563670225644, 0.0189527728602388, 0.0128785991437561, 
    -0.150062520037214, 0.0724524646348775, -0.113928920318629, 
    0.0147655867538117, -0.0134259545048549, 0.103388241018739, 
    -0.17944413876531, 0.16514602292943, -0.159453617835476, 
    0.163369165108908, -0.0309103671240678, -0.000139344881472478, 
    0.113600510327041, 0.502621995374437, 0.204751188218202, 
    -0.27052867241161, 0.322206505900714, 0.380762743432688, 
    -0.288952081530039, 0.321652421614055, 0.642337805261031, 
    -0.0661279267800443, -0.217027595097338, -0.110772442955674, 
    0.546157475643344, 0.00368459687546394, 0.819025835027298, 
    1.01570189085137, 0.0493300081483758,
  0.42748525314986, 0.537545872335194, -0.193887315595194, 0.414217026687727, 
    0.767404648359344, 0.123626223981417, -0.290389445934572, 
    0.0930331699560484, 0.581305630661338, 0.327104785234226, 
    0.409390028803749, 0.596930236950853, 0.23164703723606, 
    0.0868085334867321, 0.0222381288240232, -0.0296007469767587, 
    -0.0491315732101705, 0.516654395494937, 0.256164451250884, 
    0.0134512155611588, 0.213408915506533, 0.235837473600549, 
    0.174034578936008, 0.407666828743522, 0.159448661702219, 
    -0.07947845222864, -0.0615447803925734, 0.487085476584589, 
    0.0556260905274844, -0.0567503613204393, 0.106792304076206, 
    0.119376872706677, 0.135052902159787, 0.410698834168195, 
    0.131946008235828, -0.0685880288127339, 0.0154110977067397, 
    0.336255981600003, 0.0329287281764922, -0.0932138270243265, 
    -0.0601418881437908, -0.259278011351441, 0.102843951980963, 
    -0.123014811970055, 0.108218067738453, -0.148903049196143, 
    0.126771011007945, -0.10632056607996, 0.108602933099152, 
    -0.325040253055695, -0.00735091144790603, 0.0100901683537969, 
    0.0299258495683195, 0.0972623772775136, 0.127539302504978, 
    0.0694327167319836, 0.0149972457804749, 0.105295305344796, 
    0.236875451778941, 0.124912952193319, 0.0617977761607276, 
    0.361248969944233, 0.218900795035533, -0.380076100908403, 
    0.21016059888393, 0.947642938689901, 0.0911966804947057, 
    -0.189123508653687, -0.0647231964338805, 0.182636141533285, 
    0.893480623091153, 0.421988465311079, -0.144193880446377, 
    0.0991597866361269, 0.728415750603151, 0.663278068726458, 
    0.11415210561208, -0.24345390869581, -0.0556743081630829, 
    0.657986892365313, 0.0938843442913627, 0.0274646338358356, 
    0.296858017611732, 0.102488304817002, -0.0665353611637949, 
    0.173136378945406, 0.156624301686936, -0.14483791037301, 
    0.0229998358558559, -0.253423907145074, 0.06912266925598, 
    0.240754133189258, 0.221544028985068, 0.228789740345446, 
    0.118669509747895, -0.0189236438092715, -0.150618907521319, 
    0.166764573258273, 0.293526646957736, 0.112850659463177, 
    0.173269756107403, 0.512025231856737, 0.183527769931562, 
    -0.104939121477342, 0.267669258219033, 0.272454407343603, 
    0.0139672533360136, 0.266682412296821, 0.429616240978216, 
    0.138812886933931, -0.000742430524686907, -0.0129159490241084, 
    0.0525272158972184, 0.0413099597509323, 0.0614583658405441, 
    0.0176808455021012, 0.0355915807288016, 0.0693754087435964, 
    0.153384257201345, -0.0673913527018528, 0.382902307820079, 
    0.21017880559246, 0.0468712309566599, -0.166523486865492, 
    0.276800714355458, 0.399567655714558, 0.288119923332457, 
    0.13636546317458, -0.230972189954973, 0.124265373638442, 
    0.620453819207512, 0.248563776709613, 0.519372726636188, 
    -0.315465188293567, 0.876158115655988, 0.203432382706586, 
    -0.089296206425129, 0.0406689588450914, 0.522275718859436, 
    0.376199081426181, 0.462866169144168, 0.512653476937666, 
    0.109973192340855, 0.0136944853961982, -0.00545750121835176, 
    -0.130035748985038, 0.0265923286974679, 0.280216776019135, 
    0.121094793223248, 0.0122978924198962, -0.0759968781811692, 
    0.0236548929895225, 0.221236140463255, -0.0120948735376139, 
    -0.0700622461023529, 0.0323596655747373, 0.0955342916069564, 
    -0.015056056621534, 0.0189255010719649, 0.126194621774121, 
    0.0783468543969695, 0.0781934659460257, 0.0702295456248331, 
    0.00549903049711961, 0.0632129265937274, 0.0577685886662881, 
    0.04076441212976, 0.0585439956952739, 0.0883975938639483, 
    0.0532219543425784, -0.0576386227348109, 0.0403373837106725, 
    -0.0179152783935422, 0.0250956938407823, -0.117321474531219, 
    -0.00689503039541485, -0.042537367942017, -0.0795431875933055, 
    0.0926255554929669, -0.0927398510035582, 0.0137199704650252, 
    0.0991907829377903, 0.0938983021759647, 0.100571935115057, 
    0.159689153572927, 0.136762738352497, 0.16501175254926, 
    0.261403042625135, 0.14745644616712, 0.0249125096669528, 
    0.684816520293298, 0.132388295828096, 0.00340622209663539, 
    -0.163630967204755, 0.54526100355534, 0.3089908931995, 0.349609203799512, 
    0.299423164487863, -0.21479864237006, 0.0925790597475732, 
    0.454281441963926, 0.506293422094991, 0.220452608529883, 
    -0.148120069075762, 0.0791404268937166, 0.434592164266202, 
    0.230055797893297, 0.0200468840881165, 0.561144660490871, 
    0.0496633326328947, -0.345130513268875, -0.0281968976854939, 
    -0.238795454707209, -0.0602292549330014, -0.235654241302613, 
    -0.178339370633049, -0.111557099842398, -0.255994302527359, 
    0.144340282964682, -0.196944586907214, 0.174157762828646, 
    -0.00504193384721878, 0.137465008298313, -0.132527772277264, 
    0.0631941067867195, -0.200045335438731, -0.0660825639227719, 
    0.00577871397189019, 0.110866034795792, -0.179932772183851, 
    0.0707809827796837, -0.0237424917584654, 0.00469433611427716, 
    0.114522138822944, -0.0255546438328019, -0.0094509544643948, 
    -0.0861613604590682, 0.157828433299168, 0.0553472323713252, 
    0.104768627502318, 0.281260828027227, 0.109075054204928, 
    0.271191473772106, 0.245571513134728, -0.170062778577826, 
    1.02940117484804, 0.237546259200415, -0.0112759465822268, 
    -0.401154451437938, 0.632849068112569, 0.699861849430165, 
    0.0575742192057783, -0.115753463942414, -0.151239086368215, 
    0.547455173824303, 0.270927282682998, 0.0935331040389663, 
    -0.191536688632732, 0.0704707321570414, 0.597054567515849, 
    0.0969558253579112, -0.0966877061301183, 0.15581222894505, 
    0.342773180267021, -0.0547674823063944, -0.0498930853826022, 
    -0.100791059829526, 0.0920002945321568, 0.170911911056864, 
    0.0859199958219884, 0.0701885639292387, -0.137811086922342, 
    0.233298571864568, 0.185443778469517, 0.0522722173741014, 
    -0.00302168078198298, 0.185051728285644, 0.252595905967721, 
    -0.167304761788589, -0.135982402179113, -0.294889412907571, 
    -0.0412238230884229, -0.209249408845959, -0.191035128752972, 
    -0.0696433855857352, -0.207205134552045, -0.0366426642918935, 
    -0.178608526412174, -0.00633935335522791, -0.156713473861824, 
    0.0261121324490785, 0.0302555974485384, -0.00337153183463611, 
    0.0221798128183184, 0.0415889322791289, -0.0158811350465614, 
    0.034226121864544, 0.0629688539344379, 0.078826996642101, 
    0.0224088379812703, 0.0687862289757042, 0.0963203541599749, 
    0.144402291086265, 0.165778703151108, 0.129209643746021, 
    0.0873280513283845, 0.123485443967825, 0.201942706473951, 
    0.12939009146731, -0.000970445618052637, 0.12585655492441, 
    0.35525464958202, 0.192671882986835, -0.0626799905293929, 
    0.269662632611904, 0.473754774011655, 0.166390013714683, 
    -0.0824388173826178, 0.297562645599328, 0.503054344090414, 
    0.24675930057343, -0.271691823136591, 0.437142165387569, 
    0.671033471035276, 0.163116997644564, -0.0308716554798309, 
    0.244202012371252, -0.230561263307946, 0.406009781714742, 
    0.769432101253322, -0.0245126537472807, -0.0529197946072996, 
    -0.120841184014065, 0.147311668039518, -0.0425665120446995, 
    -0.0151666581266646, -0.0875582085105632, -0.0257137464889012, 
    0.152306995459736, -0.023290643995053, 0.0213772988825781, 
    -0.146155317302571, 0.115249267028768, -0.190830757788831, 
    0.0360282902995385, -0.273558530437335, -0.0586386431770694, 
    -0.153833053257706, -0.0591333264272495, -0.158451516052414, 
    0.168977709002831, -0.014514444234424, 0.272369759504304, 
    0.320823154767813, 0.0702229133835207, -0.144078869331784, 
    0.0142152061991423, 0.323212542006678, 0.108031504926613, 
    -0.123776872522721,
  0.0409624554759674, 0.836083110519169, 0.580037757059834, 
    0.0917742913108101, -0.116614210263051, -0.259170689464401, 
    0.770791472576906, 0.342837167492119, -0.0059505224581971, 
    0.375842990770897, 0.34162663188868, -0.0434772018862819, 
    -0.0537275233196476, -0.0344768794872659, 0.280919394327511, 
    -0.0348962323477369, -0.149162975056184, 0.128886087524056, 
    0.120269506979986, -0.11336026941333, -0.0639109685190154, 
    -0.16048487881976, -0.0394689229555062, -0.120135761596079, 
    -0.0885415758988338, -0.0663153588152162, -0.212545137597839, 
    -0.00658760843139691, -0.213451456733453, -0.0251658057719153, 
    -0.0845486277718108, -0.0233583258166877, -0.0452994033460813, 
    -0.055129739144742, 0.0305005521676303, -0.0517545326825305, 
    0.0401653268360494, -0.0154553181516403, 0.038018932631394, 
    -0.0598885245811743, -0.0278090992910599, 0.150987460786383, 
    0.128253268042536, 0.0129077948951929, 0.0929551251548257, 
    0.256413854958246, 0.212762807978268, 0.0673327529803299, 
    -0.000314761522819923, -0.0674942400645047, 0.242368552920002, 
    -0.0504764305695667, 0.857036345299108, 0.337496207628654, 
    -0.0836669503157275, -0.152213538710819, -0.470572572503449, 
    0.578985962829843, 0.834426115369631, 0.164967220757581, 
    -0.138349393884353, 0.112968512352494, 0.139701705964295, 
    0.0620458807609127, 0.49713088369163, 0.263384305354571, 
    0.0236686256509568, 0.173715771620431, 0.315148604341334, 
    0.0389231915036258, -0.0225176151626134, -0.0179067043402295, 
    0.0020755274331213, -0.0149212942462335, -0.00871810656543948, 
    -0.00370465153352671, -0.0198793852185249, -0.0132934791825717, 
    0.0228705536318558, 0.0609700243930931, 0.125883332437099, 
    0.100184809958885, -0.0376785642521287, 0.241998852989906, 
    0.280001732910507, 0.220731807847155, 0.661843634885189, 
    0.322957259795006, -0.133706982903465, 0.176988453121195, 
    0.516278238578858, 0.226830291054838, 0.157267928150167, 
    0.281868814012547, 0.304083042941501, -0.368807951423538, 
    0.50173050024883, 0.546636099052023, 0.335730949398624, 
    0.125005413646776, -0.15142499600532, -0.208563145954057, 
    0.048067671705737, -0.0250785917426162, 0.0579767333927482, 
    -0.213246627872815, 0.0238552977667182, -0.0704940910018265, 
    0.0708164277763995, -0.225553709455739, 0.019817127782624, 
    0.114208772570824, 0.36215930152108, 0.228381725897853, 
    -0.0990570573568039, 0.115584950983387, 0.651048443446853, 
    0.298750710444257, 0.0703311590330854, -0.0165308701979999, 
    0.234053246690753, 0.477173311192752, 0.419618049249826, 
    0.32789162406832, 0.291853793078629, 0.244992488794337, 
    0.183145362452716, 0.18647452292684, 0.299574010277827, 
    0.293970552146933, 0.164216276616158, 0.119679573581441, 
    0.102099055783918, 0.10511996317305, 0.133112601320725, 
    0.101312034515076, 0.0736290002133131, 0.232967426469195, 
    0.0763268283279607, 0.0056862895617731, 0.145477747690465, 
    -0.208151606617808, 0.0926890613842459, 0.42300347375644, 
    0.273520760704105, 0.411874009993119, 0.457801772545544, 
    0.0976269657673697, -0.110072454856609, 0.730744782012604, 
    0.204664650228644, 0.0370379556763235, 0.017805245909535, 
    0.0137776855421171, 0.0239550010930009, 0.0221983600635868, 
    0.0219637300876188, 0.0172348539666583, 0.00934219223185018, 
    0.00835391059114267, 0.025369230940044, -0.0249297434085466, 
    0.0425976399611219, -0.0319230808876025, 0.014020438915861, 
    -0.0129545261848662, 0.0218505956191556, 0.0045619412302422, 
    0.0486466432621896, 0.0300253599153306, 0.0399079960654783, 
    -0.0814172883932705, 0.0394898582594091, -0.000454573600015412, 
    0.0707264146410719, -0.101920496898801, 0.0521654765840965, 
    -0.0653907107573167, 0.0447110273737491, -0.049403768230105, 
    0.134526257477854, 0.0582304213101902, 0.0417584620812495, 
    0.00959777006056271, -0.0577289648389282, 0.0824118998182524, 
    0.240387764926231, 0.0908674923989041, 0.133956945993504, 
    -0.0215027201961597, 0.665029175501452, -0.039630587269911, 
    -0.19782817133005, 0.0919011982718525, 0.578556771969532, 
    -0.00762607850397858, -0.537334825970508, 0.132579397616753, 
    0.744157685640117, 0.350990721503287, 0.139739465698335, 
    0.108616938445873, -0.0578511862734599, -0.160185341972857, 
    0.559982779555181, 0.457392747555758, 0.158128664279862, 
    0.0631828020003539, 0.366977913027696, 0.441339414657874, 
    0.322694344419986, 0.345454865970249, 0.182310777581866, 
    -0.208218366271917, 0.19354575093506, 0.541467067774361, 
    -0.0875476948679934, -0.0117652398604434, -0.0150320893026381, 
    0.477365742390674, -0.0840846097757344, -0.128655063866789, 
    -0.122808462960181, 0.460848342998517, 0.43500463328549, 
    0.347188637670127, -0.200058511630028, 0.26620488814178, 
    0.31422130410676, 0.0465163467607834, -0.0595687608136118, 
    -0.292008082795317, 0.0826687701382519, -0.0758526284393118, 
    0.0586721554791454, -0.247893339774008, 0.0768515528218814, 
    -0.161499258665883, 0.0402212633401449, -0.292957032447565, 
    -0.0335111960052454, 0.0394968499245913, 0.181103567043661, 
    0.176780975923277, 0.04611022931096, 0.0392500530659782, 
    0.375597096903633, 0.321425304042708, 0.0789653919994001, 
    -0.255892606210921, 0.0420713593349273, 0.276855237546815, 
    0.490010578035788, 0.680006959212149, 0.189902164669711, 
    -0.0954269403794573, -0.264622140955218, 0.871252200785256, 
    0.244738726989172, -0.223835335570901, 0.336932957337932, 
    0.642194838586701, 0.348894368557741, 0.240200873245621, 
    -0.144615670152208, 0.624218211280444, 0.195461803303132, 
    -0.0380992784255958, 0.0840789478486371, 0.524422630797979, 
    0.076876379040959, 0.00553656699198343, 0.00281599318780595, 
    -0.132516047067512, 0.241437488613331, 0.104346005938562, 
    0.0848332664988106, -0.075431232819344, 0.203500061169943, 
    0.067852726793768, -0.0321741973292685, -0.0798385361628465, 
    0.0669359167554198, -0.0486943847574443, 0.0892991370275502, 
    0.0612209572503568, 0.00269850009622359, -0.0023546874185485, 
    -0.138236851657313, -0.0873060700701759, -0.197732988231777, 
    -0.03189958628758, -0.131910413198778, -0.128861366409418, 
    0.134850816446815, -0.18566746963555, 0.052198860834271, 
    -0.116195786416863, 0.00784427473708632, -0.182795496238522, 
    -0.0196196039329889, 0.0676087260728004, 0.0661809816383499, 
    0.11120882691059, 0.184439962492969, 0.123281926534021, 
    0.0573605100453647, 0.250341496824888, 0.267287232455491, 
    0.0410356697302448, -0.0572576578949397, -0.0828543088627049, 
    0.57840326505977, 0.28725123830819, 0.180070886400823, 
    -0.258831514296096, 0.281442803237459, 0.479309363035957, 
    0.217914325897611, 0.163031810931985, 0.670184781767955, 
    0.0265018679231006, -0.426910672244145, -0.0840078506019336, 
    0.822990269970277, 0.16944442884227, 0.0735646716515805, 
    -0.196375865917644, 0.657336773370582, 0.279921581357593, 
    -0.0280454861057336, 0.1677839643675, 0.110993784324007, 
    0.554568860535882, 0.00620773967653213, -0.299904532765413, 
    -0.425754382497362, 0.0349621585981699, 0.263016561419287, 
    -0.26193467373539, -0.0456738358449564, -0.0665009087901688, 
    -0.0837954039777751, -0.0719258893071794, -0.0722579725916617, 
    -0.0732862671522774, -0.0601309836476591, -0.0659902310173833, 
    -0.0548025489341818, -0.0296586594753791, -0.00381899938779504, 
    -0.0910270853706865, 0.242227534009479, 0.326053322242832, 
    0.106470379645485, -0.081673391930041, -0.00369736673843031, 
    0.116563705839023, 0.351746873658874, 0.161393335629791,
  0.251889573160194, 0.246899650188575, 0.242900963020918, 0.222857913207038, 
    0.21212394592942, 0.218586049814496, 0.237635181419787, 
    0.257794733213095, 0.232868870811965, 0.182263693640562, 
    0.178477692807638, 0.207113174779289, 0.269315248246217, 
    0.343670232275027, 0.20732807467919, -0.0334556254150874, 
    0.213234073645479, 0.40611999159955, 0.394272180823535, 0.32992050900476, 
    0.091286889443509, -0.152158843274492, -0.173935161088294, 
    0.68313856052974, 0.228417857493667, 0.171127114456685, 
    0.259369772679306, -0.0122237970373199, -0.192712465641659, 
    0.8723076288446, 0.219400150113871, -0.060914902520648, 
    -0.075033583705196, -0.337313492449921, 0.070785208231366, 
    0.575453308665665, 0.18853204743476, -0.0623215508628697, 
    0.292532123598774, 0.243143751523051, -0.00395645260560519, 
    0.00853656342369086, -0.0584296706562874, 0.0351311241961385, 
    0.183371144573529, 0.0973512690612878, 0.0238658930687579, 
    0.0357965889445206, 0.170037023807632, 0.146949335649224, 
    -0.215644882672901, 0.429853181369734, 0.405674625457904, 
    0.173230466764171, 0.193059695827931, 0.174607168189465, 
    -0.214652415439834, -0.103233459514275, 0.700019591009707, 
    0.23680970801166, -0.021172814615806, -0.110876497390608, 
    0.192058623319001, 0.227393548455183, 0.0123062275269883, 
    -0.0398099716259403, -0.00058159003032407, 0.126187585638305, 
    -0.07670801332518, -0.123813409531431, -0.033070912207254, 
    -0.224580004156033, 0.0409651053726496, -0.180575329740494, 
    -0.0253340273221692, -0.138400703933726, -0.00528098220815229, 
    -0.126050040390068, 0.0170709277038883, -0.2522668436383, 
    -0.0475203135398574, 0.0422447397919984, 0.0168764834585375, 
    0.0675328968529444, 0.111309354359449, 0.0243177511781287, 
    0.0821751256892192, 0.211877856226062, -0.0374889417759439, 
    -0.244743972278356, 0.0396630935803107, 0.484621064458835, 
    -0.0329755513628856, 0.0646312050951353, 0.890295174616275, 
    0.147793732054126, -0.0648713994357924, -0.137028072141525, 
    0.530788047690047, 0.495840031700221, 0.230721021420935, 
    0.195360541575154, 0.0863780857168779, 0.065643898193589, 
    0.0669289075574308, 0.0322924197241168, -0.117167007864704, 
    0.074552395195602, 0.124945364106133, 0.0241785477460664, 
    -0.0663014983701979, 0.0474095283011381, -0.0831895387109249, 
    0.0524768940437952, -0.207394241422186, -0.0112413725469147, 
    -0.18804616447093, -0.133488574553606, -0.0404094773037039, 
    -0.111300651991343, -0.109551040830787, 0.0856469079616504, 
    0.08964509944701, 0.00778925811918221, 0.109324070056719, 
    0.0466189195613472, 0.205615857458751, 0.230891493017538, 
    -0.000521971723589143, 0.233889268149779, 0.264894014496104, 
    -0.049959696784197, -0.292678874824198, 0.109036793094822, 
    0.356175654396558, 0.780498122810046, 0.275695462862704, 
    -0.20403331169406, 0.406395143119555, 0.23113916511862, 
    -0.503247397870922, -0.186577101201852, -0.0904405712283862, 
    -0.258523683173875, -0.157956209570056, -0.15046341702846, 
    -0.289982646823124, -0.0830244617649162, -0.111489417546765, 
    -0.233119563879449, 0.208418430357088, -0.132036915672558, 
    0.0725042201102363, -0.0806350641011935, 0.0943741923506961, 
    -0.26905220013407, 0.066470576336249, -0.102437951557089, 
    0.0294943640770628, -0.299347276790656, -0.0555710385120767, 
    0.031675817026717, 0.0409908717955593, 0.0756571314120621, 
    0.0926018911273126, 0.079585989696347, 0.100430164001219, 
    0.126837214322722, 0.0799272417341032, 0.0107115143536845, 
    0.116601067064305, 0.203279366860752, 0.183255818158557, 
    0.17253460242247, 0.225742491575258, 0.207185569383612, 
    0.333041900027561, 0.310414746046883, -0.0225615197114516, 
    -0.0381754378496836, -0.355827890664613, -0.114583686241202, 
    0.672642621965398, 0.323468264297613, 0.183275254785685, 
    0.512703369389498, -0.308427026786704, 0.383195246275925, 
    0.968696182448191, -0.0912957042758713, -0.11444897383444, 
    -0.153323998902868, -0.0085757121118452, 0.00166629839837701, 
    -0.0414531130860001, -0.0647318588829464, -0.0296543478696724, 
    0.0171869180191369, -0.0494281500462039, -0.0625121360105266, 
    -0.0255478097504599, -0.0197487853171628, 0.0583974577977592, 
    -0.0890278303335065, 0.0441528278789558, -0.136858902957102, 
    -0.0270020891138865, -0.0236085074082908, 0.0999748482756064, 
    -0.12747788837812, 0.111489272660402, 0.131802763116247, 
    0.0402320585440876, 0.0457326999308814, 0.179115671793168, 
    0.167491796194755, 0.107888995895399, 0.241943487196897, 
    0.263318577077447, -0.145051866016405, 0.450706058606675, 
    0.361088383503412, -0.0851228788395482, 1.25928534697549, 
    0.79665082973703, 0.473379198094661, 0.455991027233484, 
    -0.15917115742348, 0.867425849866418, 0.370030565849085, 
    -0.0503118459291108, -0.0734683983721773, -0.140527775907319, 
    0.213897925278648, 0.106461489221573, 0.0402824807467314, 
    0.0795150259491231, 0.0242996296612709, 0.0575024298977149, 
    0.286787600196544, 0.0761723950834501, 0.000564066569727031, 
    0.0153497422107572, -0.0438210075250002, 0.0594753494484169, 
    0.0697711327631621, 0.0328061574552961, 0.0119119110426403, 
    0.045185985036225, 0.0149849423625356, 0.0594352285987499, 
    0.155142003664571, 0.119862247309158, 0.0389029977159287, 
    0.242403567330537, 0.280885812287347, 0.12485692230878, 
    0.0552283931495917, 0.226227748940375, 0.22575776185471, 
    0.116177406861977, 0.077899701636941, 0.089053799918624, 
    0.111856961688986, 0.118800490318449, 0.0865673682495074, 
    0.082368644764564, 0.131342355099581, 0.118965997240435, 
    0.0689290277594552, 0.132348680114626, 0.172107099861839, 
    0.110672528286226, 0.021433140324468, 0.539935535321688, 
    0.267151010652499, 0.0458087236290485, -0.0408266499742755, 
    0.475917435047916, 0.178157155769459, 0.0305513201679824, 
    -0.0374298344409777, 0.630330153818073, 0.296904105666471, 
    -0.0212663374916844, 0.300723003291202, 0.604239730240462, 
    -0.256634754024369, -0.494800345683269, -0.129299440581731, 
    0.394678125686158, 0.163916869110539, 0.0564699977712266, 
    -0.00720092273599075, -0.0743364274012182, -0.1108396057802, 
    -0.12798670680826, -0.159437812379435, -0.0922712619067737, 
    -0.164371228943612, 0.0525600824662118, -0.0562745816116884, 
    0.0330613204911098, -0.0461663758512696, 0.050483609377581, 
    -0.0269587427796662, 0.0731362863032864, -0.00789678334810492, 
    0.0780390673951503, -0.0424964764916171, 0.0455016633992749, 
    0.0689614460895099, 0.0798256932729883, 0.0872757731905722, 
    0.0900926157875575, 0.0885075621486578, 0.102506548678658, 
    0.101100347104325, 0.0676008916192233, -0.062156191935352, 
    0.332825747498172, 0.256538866735747, 0.0909705089904426, 
    -0.174666025983314, 0.0651838104780872, 0.395858316118877, 
    0.353241027897713, 0.359028783757716, 0.210688601032482, 
    -0.1526595747391, 0.139790948547471, 0.165784143050048, 0.55262052698576, 
    0.544007562658907, 0.085398028548893, 0.00261391025049364, 
    -0.0615027926941298, 0.441430507524529, 0.168430192805038, 
    -0.295965370403734, -0.317180015649153, 0.0821414301136764, 
    -0.214275739030833, -0.0116990230875152, -0.107881585325778, 
    0.124867519024604, -0.344388921711166, 0.105419860613034, 
    -0.444246008500714, -0.171350994668681, -0.0679856889990378, 
    0.0601708368145482, 0.198932825653542, 0.21444937709104, 
    0.198672960066536, 0.147215790577941, 0.114191525856567, 
    0.195587211605015, 0.294102577918584, 0.282037705261693,
  -0.0659131547279555, -0.206182794450281, 0.0520876280917414, 
    0.213186212971614, 0.161502646101208, 0.574493675750259, 
    -0.0223447519274566, -0.104381285562719, 0.31957278421654, 
    -0.07229485795904, -0.209910200712314, -0.0953161054463877, 
    -0.133665691031501, -0.156925068902748, -0.0704133122188896, 
    -0.140529097662799, -0.06960368399055, 0.0278100766670657, 
    0.174716619763815, -0.233837364055715, 0.0681423831195188, 
    0.302743746804943, 0.146854065294133, 0.0633858204047745, 
    0.0380686260237289, -0.154977750368846, 0.294306244152262, 
    0.571618224532767, 0.308591941209123, 0.0620056565267654, 
    -0.089780015814262, -0.161241422857299, 0.4724355131985, 
    0.331742081978157, 0.109810348290298, -0.0943350355785358, 
    0.0586313618041894, 0.463714178308124, 0.388019913411855, 
    0.215720638378295, 0.153206830021456, 0.248663012697187, 
    0.289752481387259, 0.37173542814871, 0.319449605304697, 
    0.123830991012822, 0.401223342196005, 0.546272061850997, 
    0.0698191298441826, -0.0678405171979245, 0.0729488615964593, 
    -0.311370556968913, 0.402158460451641, 0.758142207104222, 
    0.136092681197945, -0.0408149542032086, -0.294617736901884, 
    -0.129182228079767, 0.894468295016945, 0.223395687940249, 
    -0.027578277466697, -0.0324324287509817, 0.0514546459990975, 
    0.171030565117677, 0.452920987139361, -0.148652410493068, 
    0.501627491168809, 0.942497835607835, -0.0582740727081861, 
    -0.0945445604479336, -0.196245381998892, -0.128995196282078, 
    -0.168432895289332, -0.0960065590714609, -0.163271316839404, 
    -0.118345234006125, -0.121883150963017, -0.141910086235355, 
    -0.0404082684757407, -0.205338448884506, -0.0872763133057566, 
    0.00170244854640993, 0.303754563977106, 0.2130449654932, 
    0.0699946899301296, 0.225783233022655, 0.240866511044496, 
    0.0911560058995903, 0.309725547560202, 0.40174222103607, 
    0.18797846607437, 0.116727690115847, 0.104452859362402, 
    0.112964053731322, 0.113737892091893, 0.105385863718867, 
    0.108757792139023, 0.113020760992437, 0.125672792628034, 
    0.112212741812478, 0.0372952323319944, 0.0149964728483589, 
    0.0278482868902113, 0.0494338159861028, 0.061313407384099, 
    0.0456697785113754, 0.0700286728789818, 0.0160769620761416, 
    0.0488638429519758, -0.00176645074712196, 0.0660263817641552, 
    0.110819649819408, 0.12124655044808, 0.144400395155269, 
    0.188925744576249, 0.161554769069995, 0.113796223845352, 
    0.194376649534573, 0.26074797432234, 0.183988636801418, 
    0.129199996581537, -0.0726448638814303, 0.433574700233164, 
    0.375589293979686, 0.0964347777063724, -0.115337448869432, 
    -0.0286112589855596, 0.302081046787317, 0.599172710432548, 
    0.248662048615363, -0.175465218829738, 0.313552864973769, 
    0.366208290238058, -0.00860594865292699, 0.455686309921965, 
    0.328152113494642, -0.252338426248646, -0.0776601271965641, 
    -0.294127620475079, 0.606018442601401, 0.0684789112026448, 
    0.0182145530530636, 0.0565321060881951, -0.0967132617458989, 
    -0.0748566229601001, -0.0103099389981561, -0.0400766731804921, 
    -0.0587628439091811, -0.0173284077090506, 0.044241011539836, 
    -0.252243276899268, 0.100431693464809, 0.0219490589820717, 
    0.116632705437952, -0.331414996020645, 0.0463542250323178, 
    -0.146626982171624, -0.0533458185691113, 0.101449022764002, 
    -0.393504126573521, -0.0985989236246915, 0.0283018768478121, 
    -0.0198452066998243, 0.0952421355992113, 0.0611379022375158, 
    -0.0791416553255017, 0.00873366189251919, 0.213917401353466, 
    0.0730134610030866, -0.400890652757125, 0.129722547595932, 
    0.547678707115673, 0.136447368057851, 0.381186026992351, 
    0.355908003009246, 0.321094716056862, 0.987997245555293, 
    0.243404909604499, -0.150168523171464, 0.0915690264853413, 
    -0.443674449066137, -0.0862999266030653, 0.662769518601331, 
    0.299542540447668, -0.0722911733901294, 0.191616075328264, 
    0.446587647486321, 0.486303980840877, 0.37943865396676, 0.18626672988901, 
    0.17223345406254, 0.32718703441452, -0.113905138616488, 
    -0.142178275112823, 0.0218473744017143, 0.0767425968051366, 
    -0.112696869857969, -0.159371395529241, 0.0417435634018841, 
    -0.0512364514201871, -0.105818327139642, 0.178331312534181, 
    0.224806331717373, 0.186319469676036, 0.128161613676798, 
    0.0422348656210632, 0.0972812433192764, 0.133241322662274, 
    0.135301024894245, 0.0494195191457871, -0.0491378098963214, 
    -0.000852227859850035, -0.0405303169902638, 0.0296669831667564, 
    -0.0433873169425486, 0.0246226007952889, -0.0247579140824109, 
    0.041854760776505, -0.0759056801682781, -0.00720825713664702, 
    0.0212650132169669, 0.0681613452722836, 0.0578255836800861, 
    0.073387602844104, 0.0541434827544492, 0.0682296661254821, 
    0.0419271479995887, 0.0569655081380151, 0.0358098611864315, 
    0.00318083358062202, 0.0743117524771306, 0.114804999918931, 
    0.113687633441218, 0.158983456969762, 0.220842899334432, 
    0.167945204491414, 0.11606717327808, 0.193358417741399, 
    0.164039412951834, 0.0934699522665474, 0.498312179223209, 
    0.251842029969776, -0.149828993070853, 0.0881632793666576, 
    0.518326214650205, 0.293365801575644, 0.260212865281043, 
    -0.195854826956273, 0.298399242084413, 0.40155551327105, 
    0.241192502701796, 0.106764843970444, -0.162967800537508, 
    0.254468061657531, 0.317394703055571, -0.429325000041885, 
    -0.336548407539308, 0.00214191643954692, 0.459572419250724, 
    -0.162608250960109, -0.0728726825750075, -0.183140244421547, 
    -0.0584885704403692, -0.182052339693459, -0.118077387846198, 
    -0.192940403401181, -0.135661497591508, -0.124878350942228, 
    -0.100779077956215, -0.132496226070381, -0.0309700157831737, 
    0.0457440678510683, 0.0348300248242236, 0.0552598826488297, 
    -0.00941916563006379, 0.042317019538575, -0.016691500378041, 
    0.00644814476223282, 0.0256795023662114, -0.0299265281817756, 
    0.152130773627794, 0.190426218868365, 0.144894334758467, 
    0.012806273210088, 0.00994659798047542, 0.364002745066414, 
    0.388503753016611, 0.206178644821944, -0.0728444208319333, 
    0.484123185408295, 0.653112455870863, -0.164974360959901, 
    0.291359372663287, 0.708919237965411, 0.0735365639880608, 
    0.0982558614132188, -0.0992143488890385, 0.34091930848639, 
    0.677223906116462, -0.0692862780699233, -0.154592306515871, 
    -0.133708066557414, -0.0646587222060892, -0.112472350206256, 
    -0.0671403451175126, -0.148644353490538, -0.0991994825128053, 
    -0.126395824609808, -0.0817240679093727, -0.119697349359567, 
    0.0458330367085581, 0.112553469524456, 0.118786575280269, 
    0.098737790009239, 0.102668697638884, 0.098978787572392, 
    0.115403663221712, 0.0795050572097697, 0.0809104039612701, 
    0.069892839343477, -0.0452979680271844, 0.00870618080448929, 
    0.00631087580637298, 0.00363134118999545, 0.0871018504119961, 
    -0.0302476734559848, 0.0327818243072636, 0.0223108484106552, 
    0.0503218564898277, -0.0554591951040698, 0.00998571642897791, 
    0.145290974542883, 0.166041394163018, 0.131622774643761, 
    0.124063237392325, 0.0844904171852945, 0.119658988929871, 
    0.340920482784426, 0.33812793280126, 0.12918808905518, 
    -0.215415881664867, 0.217866835385926, 0.599501814791087, 
    0.0237080715684946, -0.209269778739533, -0.155952417913554, 
    0.675298286945008, 0.300244060225235, -0.0830947398264322, 
    0.602288838302348, 0.572894778037542, 0.146231130041826, 
    -0.0292820380175372, 0.227283019005122, 0.0976623062668084, 
    0.37119910866496, -0.331215253079029, 1.22636758721083, 0.66728649514799, 
    -0.0633983983043706,
  0.160466348959694, -0.082500225451735, 0.107235712968852, 0.35202938630433, 
    0.261836163132346, 0.196182497337187, 0.107332066047856, 
    -0.0843316409631039, -0.180854178703908, 0.602602232925596, 
    0.287811077812305, -0.0152858538744601, -0.180808818012019, 
    -0.0607968676139031, 0.982166247873067, 0.097224862853213, 
    -0.214090164475451, 0.514001436504876, 0.0381661582876309, 
    -0.258419956295526, -0.265297112665585, 0.0528210302682745, 
    -0.174064451783332, -0.00182820851881554, -0.160366121087547, 
    -0.0391277247602964, -0.19724037621273, -0.147596445700552, 
    -0.0517660229863113, -0.158989303114113, 0.0162427460534896, 
    0.0773481083267516, 0.0781406852250199, 0.0884622044389076, 
    0.0934372083018967, 0.0898949666844426, 0.0956852655579906, 
    0.0855843757939183, 0.0755547962867722, 0.0520850995021069, 
    -0.0232816285264623, -0.0769517626363681, 0.0443052196958282, 
    -0.0450140613365705, 0.0431714221151598, -0.0628824536814459, 
    0.0129990164989354, 0.000650024471180469, 0.0655097542252328, 
    0.0167395966342262, 0.210953483140956, 0.0553953999729843, 
    -0.0705656235553359, 0.153162425169738, 0.293798737110165, 
    0.148682785693609, 0.124754253913059, 0.312422857148193, 
    0.044790920243502, 0.0246228532296723, 0.579279462316037, 
    0.0772289449056585, 0.779963387276288, 0.55374939433506, 
    0.325900715457913, 0.292660040733002, -0.133569565281794, 
    0.13088417180761, 1.12782250159784, 0.20645741827529, 
    -0.0402204016844024, 0.103800905279653, 0.187961625574228, 
    -0.421021139485971, 0.401834821702507, 0.224941833100348, 
    0.0195384747807001, -0.0725750647696759, 0.395047899381776, 
    0.304154637611741, -0.0431026422946365, -0.0907221059925556, 
    -0.0594493009433105, -0.124919962269864, 0.0064355106266034, 
    -0.015291454122516, 0.0112389207746217, -0.0818317058013204, 
    -0.0537237674168414, -0.116063871074971, -0.0108857727495262, 
    0.0587795873864461, 0.115843528052126, 0.20752835099786, 
    0.194954334201076, 0.0933192315574756, 0.108210491244405, 
    0.280712625494259, 0.14164411081979, -0.0925498898598033, 
    0.436393819813611, 0.290680656737294, -0.0836311440018642, 
    -0.165585145916366, 0.547883046943126, 0.35869245708065, 
    0.179384217922824, 0.114984656356078, -0.211012641854138, 
    0.585179379308438, 0.209201033234228, -0.0267477748560211, 
    0.373364243730782, 0.42093199492564, -0.283174067948182, 
    0.314233595447504, 0.731230008923356, 0.000589715614899122, 
    -0.1985520987381, 0.040941292593171, 0.401737714233331, 
    0.242512502523478, 0.110495337078802, 0.110871472800072, 
    0.218185576747514, 0.140912159282948, 0.0258685051328478, 
    0.0912804649947313, 0.216844690521928, 0.216952996382575, 
    0.163766724394568, 0.0259600587761937, -0.215563441646559, 
    0.379233492146802, 0.417868722035215, 0.140824743795656, 
    -0.129500383454462, -0.0187647047360456, 0.312960106383122, 
    0.406074481468889, 0.336643597284119, 0.0900421521460641, 
    -0.163291904429701, -0.135556420720351, 0.216527896430047, 
    0.425104106465788, 0.40071989533319, 0.2095460513595, 0.214264448014029, 
    0.582804571646276, 0.0358173985057884, -0.0264476053468217, 
    -0.0270351405907363, -0.0242767394256744, -0.0248322469704918, 
    -0.0239387956378424, -0.0229825277011416, -0.0212749007855862, 
    0.00400707478051401, -0.0293819078184963, 0.30367757804986, 
    0.0685365867945885, -0.0862090181617482, 0.392981417622611, 
    0.363091438794465, 0.166672670405307, 0.068969380950344, 
    -0.17477610058448, -0.0106660800741845, 0.538780110331665, 
    0.217887203247052, -0.0539693225910842, 0.0384034525713333, 
    0.311231436611347, 0.49570638863742, 0.273880613163337, 
    0.00839432094258075, -0.0105726789868414, 0.722235116835615, 
    0.135537232545724, -0.0252598747299019, 0.0328367106013897, 
    -0.0602895549528168, -0.00423006005082553, -0.00433241796739935, 
    -0.048276178593211, -0.0215350742295727, 0.082416325708659, 
    0.104465654523042, -0.16007362360258, 0.156114381527007, 
    0.325414639573095, -0.0321109667555516, -0.000643088429687813, 
    0.462412066545118, 0.398663825526453, 0.23884932350086, 
    0.0474598371829327, 0.552297430416903, 0.131788664816637, 
    -0.0612636334376223, -0.0293234847257783, 0.0526519148969613, 
    -0.0658783125371753, 0.0166625305187024, -0.0360964030505003, 
    0.0216589467459544, -0.0482805436965914, 0.030756010696649, 
    -0.0568792246295757, 0.0272026981964244, -0.0727195498139523, 
    -0.0143179557470421, -0.0284496713973654, -0.0407132676902968, 
    0.00145058197365622, 0.0406191127726695, -0.021355290993487, 
    -0.161429924771395, -0.00197551637490435, -0.284215003353514, 
    0.352595421863752, 0.407339776657426, 0.0773234942636485, 
    -0.0250285027531735, 0.365886844863523, 0.0491386289854048, 
    0.840091815475836, 0.079754543022769, -0.145067967422225, 
    -0.183227532754485, -0.305918408067492, 0.787568813234869, 
    0.797661669825583, 0.203881010105926, -0.675237598650441, 
    0.421485682591612, 1.02484274823335, 0.512600945200432, 
    0.677239510147127, 0.664222185122804, -0.146283664926546, 
    -0.0613576246571515, -0.0822574967315648, 0.000184497216800958, 
    -0.164886555428553, -0.0103784916928642, -0.0176428405177755, 
    -0.0144050075170852, -0.194403484611318, 0.193149105980784, 
    0.233372624261997, -0.0988061080203207, 0.217362202855566, 
    0.414967171489482, 0.112793262191417, -0.0155401545944036, 
    -0.113796280607962, 0.17028254240603, 0.461285199237084, 
    0.270038167800903, 0.0366317238318882, 0.0976177496412871, 
    -0.0287455450848546, 0.228263600831769, 0.939335740820929, 
    0.201901039901874, -0.234685402011242, 0.0945470305209442, 
    0.746934895985804, 0.114801643919645, -0.134735676779125, 
    0.342329439836001, 0.299832893554367, 0.0284940929548942, 
    0.21035198004541, 0.344081202805837, 0.80711400599222, 0.327064332725763, 
    -0.173870656561768, -0.13886620569815, -0.129903615931336, 
    -0.0553176712684525, 0.0844094680706774, -0.0355105374104509, 
    0.169790958815078, 0.0836985871111238, 0.00413277194875113, 
    0.144001944450344, 0.0833611873750063, 0.0347449667679204, 
    0.0338583731720314, 0.0280681725712586, 0.0337723430209315, 
    0.031183663206804, 0.0307130902504197, 0.0173596591446151, 
    0.0583092708774628, 0.135916497723601, -0.0700506597389298, 
    0.475059219853187, 0.120354101368606, -0.16175274284744, 
    -0.00993120979837693, 0.593066717407885, 0.108968037456914, 
    0.0131787720532915, -0.0688538740313063, -0.197699411409535, 
    0.380161677058297, 0.614008299726132, 0.0887050866976253, 
    -0.0556535476197297, -0.0146562003078713, -0.396189280882037, 
    0.73773469572551, 0.415808108798194, -0.0240871218515706, 
    0.511980422307313, 0.476035233053239, -0.023191830978206, 
    -0.0639501956679513, -0.0637470949825995, 0.418377934067045, 
    0.146548234515481, -0.0351546140438692, -0.0159174476475678, 
    0.307133245120412, 0.219594585440865, 0.235604112627414, 
    0.34005994208164, 0.185743030303143, 0.266739603857031, 
    0.230408561791128, -0.131962550135173, 0.196597712872602, 
    0.237334876395258, 0.0464217632342167, 0.262807636990065, 
    0.301193024078756, 0.116531293714129, 0.0741250693975404, 
    0.0319605404051743, 0.00869418240011459, 0.144954405722264, 
    0.0520477236382818, 0.00617876165784617, 0.0480466916351326, 
    0.174228766772094, 0.0542217818913132, 0.0135670072347522, 
    -0.0139676157436169, 0.0399707470269577, 0.00240795959419406, 
    0.0136102024688403, 0.00981173735923069, -0.0209043000474561, 
    0.0378595378666872, 0.020718378500224, 0.0646765310986687,
  0.0637476270432383, -0.18782344607691, 0.426666159823886, 
    0.218803967365735, 0.315244084828189, 0.887440083826751, 
    0.31645004334226, 0.129733528226365, -0.194105784690086, 0.3796149784839, 
    0.429886893529553, 0.312608030457377, 0.236425722208553, 
    0.0930634452300672, 0.0286941409257121, 0.175386888203847, 
    -0.429896388709204, 0.543542382315445, 0.387678718741894, 
    -0.131268479261136, -0.245624982245162, -0.0939529590020269, 
    0.150752567357966, -0.0487773229723012, -0.0662421472495748, 
    -0.127041148691334, -0.0386782441548067, 0.0445036480694475, 
    -0.158744560478568, -0.068166097433005, -0.0350306743134648, 
    -0.0118542409481489, -0.0270880995821376, -0.0253677253664874, 
    -0.00242424224664864, -0.029638284443896, 0.0191976842716404, 
    -0.0166143127763982, 0.0665702622316812, -0.0296363023750226, 
    0.184553917537611, 0.096716596683051, 0.0497794263958247, 
    0.316159661283191, 0.182124024216068, 0.0645553425591577, 
    0.0677175308970397, 0.216516791140007, 0.0798683921118802, 
    -0.0978142041879233, -0.0556670734414634, 0.568084280286846, 
    0.608065492321543, 0.417324998447355, 0.191718538132609, 
    0.897148239666631, 1.02172991983556, -0.115596960311653, 
    -0.143263264146591, 0.0741729162114533, 0.136442269682448, 
    -0.214212148463534, 0.0646667847168289, 0.318302938487637, 
    0.207090459010386, -0.0360573672737147, 0.149932358169438, 
    0.28234896500639, 0.119245057072487, 0.0133937071348471, 
    0.165396050664792, 0.280796457255817, 0.102302354446528, 
    0.00597305811177772, 0.0262094201347108, 0.188380873291949, 
    0.121876541018814, 0.022634705893806, 0.249151063590202, 
    0.168994816344714, -0.00830590862248469, 0.153934400171825, 
    0.39713987429545, -0.0788460057755926, 0.763105375836467, 
    0.555775383045476, 0.0281429014997129, 0.855294247556956, 
    0.465664671193782, -0.196161915586353, -0.173400634167494, 
    -0.170158630206433, 0.267968074943596, 0.199822489240337, 
    0.0324130412575019, -0.212322364664824, 0.0748327808370379, 
    0.160497404320221, 0.075033397756775, 0.294285971010538, 
    -0.227584339033499, 0.245577324017, -0.133081487994211, 
    0.207404068377195, -0.166992258778089, 0.12771677613906, 
    -0.240100035499571, 0.00311705822855177, -0.496917773107345, 
    -0.147392965816662, -0.066328966542262, 0.098507988384236, 
    0.0658489885653713, 0.0666637324204491, 0.0163629164172756, 
    0.000442143960364322, 0.0279333175651708, 0.0917767412236199, 
    0.107632405448354, 0.0391024394398556, -0.0689721249373505, 
    0.18113499963114, 0.330254012056672, 0.120361353404205, 
    -0.0387556504772188, -0.00539260811627279, 0.353478131720212, 
    0.388436322177717, 0.230546262600617, -0.148767883878042, 
    0.44435827762384, 0.363027540430242, 0.0821054148548011, 
    -0.0901964321374449, -0.163569177060981, 0.278422094635132, 
    0.594826382462624, 0.406368148257642, 0.199634924655384, 
    0.157134460627395, -0.115019259331943, 0.659226784365822, 
    0.0442147382366525, -0.112157878675195, 0.0298638369335899, 
    0.549691069531224, 0.0129614307818839, -0.050916617219545, 
    -0.170934429403111, 0.372159068729786, 0.351107641248192, 
    0.10586992162953, -0.131584344980958, 0.0169199675262731, 
    0.327983093868686, 0.202534371550095, 0.0355569321830219, 
    0.411674277786414, 0.201342948880461, -0.175978904593154, 
    -0.213319992671061, 0.0279596467302563, 0.0904521320276254, 
    -0.0342626851438984, -0.0500980752551866, 0.189028562498771, 
    0.00522874776021839, -0.0950144130775596, 0.135580871816921, 
    0.0656978437643415, -0.0401993900651924, -0.106806731778292, 
    -0.314642158468958, -0.127547179472612, -0.517363606353158, 
    -0.263232942388152, 0.0579106178576711, -0.264590828426405, 
    0.0701212561163206, -0.375909155228554, -0.0476468280377032, 
    -0.0305159801512896, 0.094298620548554, 0.152516932260243, 
    0.0882577749375952, 0.0421924013453522, 0.195503689342408, 
    0.181848277185349, -0.00781551557058244, 0.188326138459201, 
    0.470162223121471, 0.0884032414841254, 0.0429718703090325, 
    0.823116853993487, 0.354421661051543, -0.0547417815570907, 
    0.790164442319122, 0.561989123222681, 0.292285044922957, 
    0.218387035691568, -0.452931685352941, 0.073594255882228, 
    0.171369194118309, 0.613771519645467, 1.13964108926839, 
    0.0817503189362218, -0.498271607485481, 0.104685820104812, 
    0.812444202746475, 0.0590341847358436, -0.00279104186946759, 
    -0.313140678654963, 0.134830467351019, 0.443744741171614, 
    0.0510375039010835, -0.301237914436283, 0.124479362705276, 
    0.310180923410714, 0.00820869280422677, -0.0493681907753139, 
    0.325647796246074, 0.319613776980813, 0.25085695034579, 
    0.0820118758354975, -0.131564401486235, -0.150360634813896, 
    0.383298336951369, 0.288636698979949, 0.149086606623759, 
    -0.204106302349606, 0.130649608878285, 0.262108580174152, 
    -0.00141649071904541, -0.00116046669401608, 0.017461968559128, 
    -0.0608798231340678, 0.414259575529742, -0.109245468400469, 
    -0.177269907764254, -0.0100371731230524, -0.293078362059429, 
    -0.180603010238513, 0.0915334750778829, -0.120965026079689, 
    0.222070372473596, -0.147684363531075, 0.0755401897744816, 
    0.00386934423003522, 0.12657985933729, -0.20608883009588, 
    0.0479594732382237, 0.0934927524393343, 0.113461867893481, 
    0.0902252058496558, 0.0953845635756315, 0.0751184858169735, 
    0.0994426832456738, 0.158093791476314, 0.138138564145846, 
    0.0690407263113468, 0.110564847019688, 0.180201549944012, 
    0.166977247755789, 0.129585959696089, 0.198933207756703, 
    0.179472376582972, 0.0203753774383811, 0.508884706588747, 
    0.226209451171607, -0.206068647869879, -0.0575986397213104, 
    0.540655292189802, 0.501921431883181, 0.347185109167098, 
    -0.265679101530562, 0.662179266925389, 0.357240911711451, 
    -0.239901749725555, 0.610664489453361, 0.319857327995229, 
    -0.358756300973414, -0.0192437088459421, -0.147168418336288, 
    0.0114454638536085, -0.181754687215498, 0.0270484317031518, 
    -0.260197207989951, 0.144651129220872, 0.00402689340928177, 
    -0.0514831837576304, 0.0178871961414443, -0.342989200519581, 
    0.215164428288085, -0.234608902123629, 0.0827500872340182, 
    -0.317258187751631, 0.0463985281875137, -0.240836417381212, 
    0.00797828310217916, -0.398394688801641, -0.146508688687024, 
    0.11965710075438, -0.0389539845746402, 0.0907353870743898, 
    0.253296227930175, 0.0179976103438364, -0.0443744830569887, 
    -0.0926194710450981, 0.440722306572819, 0.0179972584569978, 
    -0.0519637040233732, 0.0126639198487877, 0.743850664810197, 
    -0.0259265978487136, -0.0823828152337494, -0.162879607105665, 
    0.76189643659093, 0.134629427657295, -0.0294326109334659, 
    0.0857490961485775, 0.394684728220479, 0.141433935385664, 
    0.146610063812319, 0.195703085763275, -0.122941617932594, 
    0.213995085312506, 0.279827307560254, 0.242673684365169, 
    -0.0378428324480483, -0.240334562442866, -0.283679297943864, 
    -0.0864453986351257, -0.16427153721469, -0.190227612896985, 
    -0.10707227128697, -0.157250380124684, -0.125460810016084, 
    -0.0775197525263401, -0.188696175863669, 0.042443985054377, 
    -0.160178083914416, -0.0301438931719911, -0.0247337531162839, 
    -0.126766391199379, 0.147524109223703, -0.0637682297585814, 
    0.0375471912304803, -0.16528658796218, -0.0350130838783821, 
    -0.0648526384656471, 0.0317773455537211, -0.0287259576322161, 
    0.219231175340184, 0.172482253068331, 0.0551862073532566, 
    -0.0498880426523278, -0.071709379542325, 0.183819748807357, 
    0.34621762588085, 0.113821087404293,
  0.376002733850525, 0.0353906534183631, -0.150568254920984, 
    0.533762705433038, 0.550453350163605, 0.363034754921089, 
    0.227162006613822, -0.438895574675443, 0.306544423147309, 
    0.543523971668232, -0.0443551724833883, -0.137585909173702, 
    -0.178021696158349, -0.0984289261156738, 0.539273497494051, 
    0.373621758716032, 0.503189855490462, 0.435126724111505, 
    -0.339387771453704, -0.233820622413851, -0.144602210406102, 
    -0.207396631303473, -0.0323743458598459, -0.225583828866039, 
    -0.0226026938125258, -0.28121135095609, -0.0937325547393225, 
    -0.21363978434911, -0.140970329057001, -0.102547671754089, 
    -0.0171378137479707, 0.0889083664674311, 0.0363044289624548, 
    0.0934611685585968, 0.0418234125384471, 0.0902188337617456, 
    0.0281508664662375, 0.0703551416280239, 0.0594923828764997, 
    0.0730745178514683, -0.0237192333627349, 0.0477311261017113, 
    -0.0985478472873112, 0.0473906710443732, -0.0537698242877778, 
    0.0401997578216557, -0.139076056129634, 0.0124038201429865, 
    -0.10806473528416, -0.0755371912455839, -0.00514673748703919, 
    0.0565195414746549, 0.0971545378485907, 0.135849783499147, 
    0.111330912625822, 0.010719100890674, 0.0636704377946705, 
    0.25518851500313, 0.227407103426456, 0.208689604686648, 
    -0.247515093044298, 0.147193646760139, 0.488385867707844, 
    0.227583617276909, 0.123738768161488, -0.330135175127372, 
    0.0525434413279976, 0.555847858435452, 0.223104878640766, 
    0.0425328498707137, 0.00794002309375877, -0.0868790135038233, 
    0.534919044637315, 0.302853488272532, -0.133672573168584, 
    0.52687827077648, 0.530391879451832, 0.21674200062896, 0.600045130796599, 
    0.384328269504545, -0.225661757604323, -0.126984286102512, 
    -0.0796596871290309, -0.137557795728083, -0.198837330531898, 
    -0.226655433253319, -0.118052293408993, -0.182065911242913, 
    -0.178836046439183, -0.0122459411932666, -0.13177907767117, 
    -0.0159154054102797, -0.0987722003928447, -0.12069477825297, 
    0.0916880550037664, -0.050684175830537, 0.0427423605884879, 
    -0.131741100190861, -0.0605218378180798, 0.0641679081677963, 
    -0.0758896572601604, 0.152232583226804, 0.189985256235703, 
    0.0363046688094549, -0.0212549369030103, -0.00701608386607043, 
    0.427815760654714, 0.153026912567101, -0.00526780038311446, 
    0.0213091962803583, 0.171082478978271, 0.0612284605217502, 
    -0.292064150806941, -0.0590513324905054, 0.688274893553879, 
    0.483781337123244, 0.0879663440900862, 0.392334100895921, 
    0.944022952245562, 0.14838384180182, 0.0496356530951023, 
    -0.101872466735974, 0.378345985321412, 0.234637395583847, 
    0.0965308553145134, -0.0305237130071208, -0.128658283364428, 
    0.388974337595016, 0.235876741570161, 0.0397537245010625, 
    0.0685630473817889, 0.278385674640488, 0.143075592583308, 
    0.0647657721244498, 0.0531609368353165, -0.0842671158463622, 
    0.138422554919703, 0.117780841710056, 0.0743689462113693, 
    0.425845705243229, 0.20359183478191, 0.00639273703712769, 
    0.22326532911963, 0.203731936410875, 0.0636116714760731, 
    0.116094994152442, 0.22009333113626, 0.224604762457274, 
    -0.155845631328299, -0.0853321837435971, -0.21716557059558, 
    -0.203621168376708, 0.132892544637328, -0.186675150530792, 
    0.0976730182413357, -0.137705447297408, 0.0054415980829602, 
    -0.0535528964552665, 0.0845098702524862, -0.241591168201796, 
    0.0731794367369579, -0.00120211288355571, 0.0161608464434693, 
    0.0438454815231909, 0.0579872747573865, -0.00586037475010447, 
    0.0392881178934109, 0.0303440371355963, 0.0246141891101295, 
    -0.0515405473567354, 0.00131181174170679, 0.0924586099119074, 
    0.117872058912466, 0.10057276658308, 0.10180392244929, 
    0.0891828842680211, 0.14491147509537, 0.260390599250434, 
    0.133889026494796, -0.108515210908363, 0.115928395296629, 
    0.531165629877292, 0.176449855993342, -0.237717755717451, 
    0.207617972814628, 0.504397783281197, 0.18107046021988, 
    0.0405934587463655, -0.14586775633425, -0.215134782777342, 
    0.725934462535562, 0.151394312861644, -0.0673896320887337, 
    0.00249507902813915, -0.132374927879466, 0.759241082461658, 
    0.528947462330312, 0.140716451629981, 0.709595891019468, 
    0.56610117997372, 0.156195310196912, 0.181599367282234, 
    0.165724427340222, 0.178097175318475, 0.491551954875551, 
    -0.0241990138844457, -0.221512219055783, 0.00522873055964529, 
    -0.0158302736476509, 0.339638124392634, -0.0296887934832931, 
    -0.0113008139260548, -0.0546051278332534, 0.000141020864521044, 
    -0.0485985511566411, -0.0185206546852765, -0.0388818245371471, 
    0.0579101773223537, 0.271423929256478, -0.226753649450275, 
    0.303010413858577, 0.455644901911258, 0.159677784041085, 
    0.00994056899287307, -0.16154731580562, -0.222929369526485, 
    0.373191009396193, 0.489510849179166, 0.254755074695574, 
    0.119462404492305, -0.178138319228971, 0.292208805962355, 
    0.308442949750723, 0.138583862728769, 0.137796491712307, 
    0.303836308646027, 0.0102931028714777, 0.169903085408681, 
    0.582615726404351, 0.0728586257029403, -0.0685849458680191, 
    -0.0342645199056833, -0.0285005673592891, -0.0368362720269204, 
    -0.0310901518618708, -0.0364518053218104, -0.0288443965742849, 
    -0.0289854423109484, 0.00953271662487983, -0.0837463260173339, 
    0.0636132181448216, 0.116252795013216, 0.06279618988766, 
    0.215111572794889, 0.242817850600689, 0.0731458423253492, 
    0.0766440294379741, 0.435552838225422, 0.11618779996591, 
    -0.262898436834887, 0.163828096977783, 0.586772325650864, 
    -0.00073615164746367, -0.271226288320467, -0.177548356452461, 
    0.681352518099911, 0.597728482709015, 0.165928824834466, 
    -0.149428127661342, 0.176011412282162, 0.256650216029669, 
    0.0667296067135863, -0.0154721873122796, -0.019151048452933, 
    -0.0649564932215247, 0.0391314036618172, 0.0438485029755917, 
    -0.0751070046442874, -0.0511275805879003, -0.0634953035529518, 
    0.0221585462981458, -0.0745412710673774, 0.0707318159926213, 
    -0.0836212889761973, 0.0366343461683689, -0.16261387137462, 
    0.0170427220496137, -0.0563815692721096, 0.123684909657823, 
    -0.118147561513962, 0.295170700583309, 0.132062327579439, 
    0.00464110029454201, 0.0776461658537365, 0.142459723083538, 
    0.243521839117816, 0.45017836758712, 0.421946498628366, 
    -0.00542483042703665, -0.284735529743287, -0.368123455904465, 
    0.546367602224829, 0.578500763554085, 0.211596777903571, 
    -0.398788439931616, 0.393848544406303, 0.544669877782758, 
    -0.0972840249491299, 0.287442482864544, 0.927186678079619, 
    0.441893908553392, 0.126824876750691, -0.136400246638543, 
    0.125950675093467, 0.211385169677146, 0.192783762252281, 
    0.17821151202947, -0.0676570606896908, 0.393857873552319, 
    0.149707444677536, -0.0317019921132409, -0.0256714009079371, 
    0.185039905845877, 0.162237473797728, 0.0361019988513724, 
    -0.186032312017621, 0.0528883055502907, 0.2038691538259, 
    -0.0717744123140415, 0.0133588617493568, -0.219234430472429, 
    -0.0783851046998134, -0.140567824832449, -0.098055676977274, 
    -0.125316593553098, -0.0673964873718867, -0.119687059290422, 
    -0.0229447526378835, -0.0850068660482568, 0.0171425062808989, 
    -0.178515650609541, -0.047710862136563, -0.0185796288172697, 
    0.0344053599507568, -0.126837763337944, 0.0401027107314381, 
    -0.112786703139926, -0.0560054463328521, 0.0826972195067878, 
    -0.223613853580412, -0.0184038517628962, -0.0109554729475369, 
    -0.0175866192752157, 0.00599662937796933, 0.0124841685593179, 
    -0.0209416707753005, 0.0244103687584476, 0.0288633162530993, 
    0.0411573620317955, -0.0461778119839044,
  0.474922695749893, 0.288424098251758, 0.170301012707609, 0.15727970066906, 
    0.148552106093554, 0.0869902423279085, 0.104282439688326, 
    0.247905973881074, 0.0883977122464554, -0.0629276427605589, 
    -0.0420842974190354, 0.448715589088535, 0.181943980575553, 
    0.0573270196141266, -0.148788592722235, 0.308855426710512, 
    0.304914212989718, 0.100624422163197, 0.602385221553728, 
    0.430288305384276, -0.103418734335366, 0.599401559896315, 
    0.359964300039187, -0.233253068968312, -0.280909489647932, 
    0.304631536919721, -0.478689309337876, 0.865918893193594, 
    0.567754222035016, 0.0786018981531435, -0.0234216577795871, 
    -0.313089243615445, 0.039544946936646, -0.0801150344151477, 
    -0.0882890342672431, -0.0779128149196503, -0.0392594777070862, 
    -0.0165476491121788, 0.09524120400844, -0.0316778509221207, 
    0.0107824253698838, 0.034262612439779, 0.0325893591646306, 
    0.0329221932969437, 0.0334301051622555, 0.0326463828406632, 
    0.0356541195061915, 0.0266945854639498, 0.0278481418552602, 
    0.0501564032372923, 0.226310260942239, -0.0632649814817553, 
    0.113807262786119, -0.378080505187007, 0.650505602410073, 
    0.496236372679105, 0.162811080656704, 0.104897709184044, 
    -0.205496095430267, 0.0827961626443286, 0.629615752782859, 
    0.0631475215678082, 0.0264309353376506, -0.141990129413601, 
    0.524155987760746, 0.0923264212657661, -0.144561225977633, 
    0.221691668105687, 0.318150509113163, -0.0105979090148184, 
    -0.0617791473040305, -0.162790241984428, 0.0163315161173036, 
    -0.102157396707734, 0.0152229706720972, -0.122423737382342, 
    0.035307900746958, -0.0616558167617117, 0.146751275767191, 
    -0.115365379136031, 0.417494376114156, 0.13604517720864, 
    -0.00454505959218712, -0.143127121905671, 0.127338282277359, 
    0.477497882944607, 0.419031184317804, 0.0739725668340191, 
    -0.120347310646569, -0.170641911542623, 0.207964668920782, 
    0.364321580041974, 0.789142688984194, 0.237267601563065, 
    -0.165467519440488, -0.266619813208163, 1.19287198348509, 
    0.0941641678126221, -0.37959470797499, 0.580687210419048, 
    0.405696917397533, -0.0496746854891397, -0.0528178914923579, 
    -0.113783603350412, 0.0145865392397889, 0.17831486684648, 
    0.471424660656489, 0.264596544986995, -0.0128691363093404, 
    0.361012465546753, 0.363277230319893, 0.167723644932115, 
    0.0975040923789114, -0.224186168150034, 0.137729752757649, 
    0.356418883086753, -0.0508694667079238, -0.224366662651355, 
    0.177172810124686, 0.130874781974989, -0.178118571238161, 
    -0.0289624460602671, -0.0247061706843227, -0.124544631143154, 
    -0.0280429184864803, 0.0654449458462403, -0.0122099376642754, 
    -0.0896848877497967, -0.0806434792488522, -0.0234796291336825, 
    0.0367588488996769, -0.146217246616166, 0.0820071326279443, 
    -0.0911892123117564, 0.0478810357140503, -0.124687168960161, 
    0.058427726746526, -0.0737502649638189, 0.0339639976635746, 
    -0.293404166277101, -0.0442960567543193, 0.0160258577192941, 
    -0.0107317064988572, 0.0652344332357388, 0.077665055961052, 
    0.0150026146343195, -0.0233946659979899, -0.00254472966809625, 
    0.212847559474087, 0.0683601924059, -0.109129870375356, 
    0.177978201078423, 0.587803018071926, 0.0946886281143564, 
    0.0331930125208937, 0.130598631064552, -0.490392977690813, 
    0.595971674158125, 0.567077488316772, 0.297810404668438, 
    0.599873637181799, 0.439012548527486, 0.0384736158821319, 
    -0.067752408578095, -0.245598321319042, 0.178022384817417, 
    0.550093200907306, 0.250478219164932, 0.140100250792854, 
    0.298047888207968, -0.152739075713547, -0.266196003377393, 
    -0.1497931484084, -0.204831650517187, -0.0848911305300638, 
    -0.199080620070868, -0.0032114234726095, -0.185614370501797, 
    0.0362292612933101, -0.242193451763096, 0.0444502410039232, 
    -0.00704331899199895, 0.0620479703598721, 0.0237339246251028, 
    0.0686688881801452, -0.0180734192811827, 0.0305271777999869, 
    -0.00586587096299694, -0.00159173590679046, -0.000201762059142213, 
    -0.0235311864513999, -0.073912790563964, -0.00502493431863517, 
    -0.0367160279500903, 0.0128450483371233, -0.0608160875687275, 
    0.0151040061988498, -0.0428015801909541, 0.0197210019506254, 
    -0.0792482886108931, 0.0202931418253698, 0.0557102487954311, 
    0.0864154751099589, 0.1190597817803, 0.128477723875646, 
    0.100466401896193, 0.108099342711285, 0.178609132425688, 
    0.119803541669413, -0.0175262843449194, 0.18390818205567, 
    0.300364590083132, 0.107022495478523, 0.0643142797549581, 
    0.554277366130532, 0.201363195493482, -0.0714817197309409, 
    0.0708311606527853, 0.529276589572062, 0.166954073382697, 
    0.0876192778941108, -0.0786852616593925, 0.0435328279713088, 
    0.142705960020353, 0.666936002246777, 0.420071704770839, 
    0.0664825119648832, 0.429613968992469, 0.456098114301511, 
    0.279648661212788, 0.356521076702862, 0.196420730043333, 
    -0.107255119689934, -0.120400641361823, 0.18055924273463, 
    0.083375368112109, 0.34342234092473, -0.097550790005622, 
    -0.185460521031017, -0.105705372112154, -0.069071202779541, 
    -0.268862197039435, 0.137505846685488, -0.311188966629986, 
    0.0899099161554978, -0.257969106897092, 0.0537611239123695, 
    -0.16606613978533, 0.122382846245567, -0.232463161394483, 
    0.036423042815575, 0.048646613745017, 0.055078019849836, 
    0.00410830693509604, 0.0501929839904196, -0.00344288993364908, 
    0.0348147290175489, 0.0337501303863745, 0.0545708856108237, 
    -0.041569898964137, 0.0382528270560763, 0.0890226392111975, 
    0.0787996801457547, 0.159282712200127, 0.152098395845266, 
    0.0394629014611274, 0.169546305189329, 0.259350131057087, 
    0.109174309503371, -0.0481562986029983, 0.483672696515063, 
    0.200835275869616, 0.139777687879688, -0.148090197650744, 
    0.598880055469301, 0.258264666263616, 0.416303992466743, 
    0.467612641391563, -0.102168552556376, 0.53234372332324, 
    0.322611396345764, -0.0879550215685374, -0.0502352501458649, 
    0.0550433971836932, 0.317883215632474, 0.213803883949348, 
    -0.155041361620393, 0.593930596021514, -0.20130980222437, 
    -0.223007624017644, -0.329682513347425, -0.102963861397585, 
    -0.110771775338787, -0.217916111850149, -0.0391780787075168, 
    -0.164864668242484, -0.0199212444463482, -0.226845772327965, 
    -0.0105274210004659, -0.197734632990535, -0.0720083146356377, 
    0.0733468896508668, 0.111363433792036, 0.144004355430021, 
    0.18563155117387, 0.0871090704825044, 0.0985906842452032, 
    0.394384561482819, 0.122404462675638, -0.163556522763022, 
    -0.103930464465306, 0.449257875243267, 0.70926611015881, 
    0.181024264402709, 0.0345975844241143, -0.434311246950401, 
    0.409217145936578, 0.515376711345209, 0.193693246756253, 
    0.0344162580619096, 0.6826168347783, 0.379793990667862, 
    -0.243426313189758, -0.0715576631004876, -0.209040427261549, 
    0.266460431930161, -0.133785255930357, -0.189755862765452, 
    0.378849736070184, 0.00223663554731686, -0.12864689470291, 
    0.0998211206879515, -0.356265464529046, -0.00596809106804154, 
    -0.227219302623335, -0.123313378289751, -0.125326105116611, 
    -0.0427636775343492, 0.0316538136314761, -0.234704598116281, 
    -0.101805570335523, 0.136759264345579, 0.114355558914411, 
    0.424272084735461, 0.433961407628886, 0.110428063153903, 
    0.0512306433705749, -0.352673403041705, -0.0177413750634611, 
    0.487985261630437, 0.388213520054438, 0.273306001219397, 
    0.265990344692588, 0.156305677388152, -0.291456408354672, 
    0.17449998823959, 0.672513549681359, 0.254154981877862, 
    0.00103805929366985, 0.317258263786517,
  -0.0878258800735174, 0.0391560645443559, -0.260994993845928, 
    -0.0784964454091418, -0.0179480623071267, -0.14197668866175, 
    0.076026732656033, -0.0725463361671073, 0.0745560560224901, 
    -0.162232940748458, 0.00402292534740053, 0.0600118900648095, 
    0.0446678301751879, 0.0981186393828827, 0.170767796089557, 
    0.10272248552924, 0.0462937115509186, 0.253476772420857, 
    0.178936071367393, -0.156892766737314, 0.277650854429696, 
    0.391326467389293, 0.355337508273365, 0.388430533405418, 
    -0.208226376426623, 0.594340637475556, 0.34371892953828, 
    0.0492154056527058, -0.244724326586415, 0.177683920762887, 
    0.759337254129482, 0.0708124682067897, -0.121606816239057, 
    -0.266683522089233, 0.451062007061636, 0.45391864341988, 
    0.322701998161203, 0.476180789710632, 0.351641913010366, 
    0.101087717273349, -0.19255404102016, 0.198911818743017, 
    0.412090287562436, 0.263123683170844, 0.142493066349566, 
    0.0555012199085971, 0.109558942941521, 0.231592556969822, 
    0.00331866632933458, -0.0299085767244409, -0.206897185677716, 
    0.242421459033077, 0.359054369252164, 0.155255326866463, 
    0.0283878646438321, -0.0628423551082074, -0.234506704679383, 
    0.515870081296902, 0.306540358934758, -0.0311768423615474, 
    0.469958711713912, 0.380395509945111, 0.0496245448679257, 
    -0.339974890748251, 0.0423940169312082, 0.601364899553949, 
    0.0575322652460124, -0.09227038398448, 0.178996216802638, 
    0.468750457373202, -0.232996940535381, -0.119194518285549, 
    -0.0438159338986712, 0.0392355300707011, 0.210619452631122, 
    0.0825978860041944, -0.061359935448528, 0.149706102360694, 
    -0.0589647906973629, -0.174579174188565, -0.0794994425627731, 
    -0.070035535008691, -0.084691094781692, -0.07871604828155, 
    -0.0593818739176942, -0.138964831531182, -0.028397605112325, 
    -0.114909767303992, -0.0242335561309111, -0.0633844962739941, 
    0.0348798107974568, -0.14702474528724, 0.0511802079189786, 
    -0.179365826986702, -0.049498940363177, -0.0613134329422631, 
    0.0421397491638421, -0.0902867980400108, 0.0217158716927559, 
    -0.185524715145026, -0.066987468044154, 0.0389611928688099, 
    0.0467096985922848, 0.0511479621993628, 0.0683869447587302, 
    0.0555662625352526, 0.0315303911587664, 0.0591474471134412, 
    0.044214259242315, -0.0123771691237578, 0.0827706709364281, 
    0.134070110024245, 0.137954628522494, 0.162697215260866, 
    0.189536751298001, 0.174024020731783, 0.227111961677803, 
    0.329777278405901, 0.216288842856788, -0.127845167109251, 
    0.612209756848958, 0.265250446099286, -0.0898601296736882, 
    -0.0149320855608583, 0.692773424485404, 0.265478880900724, 
    0.149388886448766, -0.238940596620932, 0.396322465423236, 
    0.630032005772509, 0.124900788458813, -0.296268338707929, 
    -0.17262104632741, 0.738728985363932, 0.214076694642425, 
    0.00549970284575624, 0.233880138051459, 0.0427546625233598, 
    -0.0107287773249716, 0.933004442628879, 0.155166841403426, 
    -0.0366266104487511, 0.0221291057837568, 0.123642707260667, 
    -0.146129242186613, -0.139923026512975, -0.0385741404240177, 
    -0.165136541842852, -0.0964621401216251, 0.0102470732552193, 
    -0.0431932136614934, 0.0173411903382773, 0.0150552643596268, 
    -0.0019525690763678, 0.0197589714107798, 0.00859828292461935, 
    0.0231480359065471, 0.0282481230632902, 0.000551207088997724, 
    0.0915435340439034, 0.25972746787871, 0.173960890619411, 
    -0.0920881288272991, 0.547509120945046, 0.281049393762721, 
    0.0566559303455499, 0.108486197148034, 0.409979591248545, 
    0.170318389822917, -0.105629684818146, 0.336685736154749, 
    0.534572559955352, 0.124034417645947, -0.0386973590843719, 
    0.117584804620086, 0.214959538947214, 0.0793228049023795, 
    0.358099661521817, 0.294236598619889, 0.00507629092816762, 
    -0.0571714529867262, -0.136383587961404, 0.0388248159642998, 
    -0.0730491375345627, 0.0268559814380376, -0.123790944155185, 
    0.0104243298406382, -0.0405299458889904, 0.0660361891133403, 
    -0.163421432240792, 0.0620233531658013, 0.114654978543511, 
    0.0171226051412642, 0.300401099545467, 0.203098152079, 
    0.0527973744406184, -0.0040742733973568, -0.0253248464541784, 
    0.0896230615275532, 0.499204465886739, 0.191472699618381, 
    -0.0402614849637837, -0.201517926999079, 0.516287538799337, 
    0.370302919960271, 0.107120328038577, 0.0364291365804003, 
    -0.25985842234682, 0.591490153101957, 0.27323637164012, 
    -0.0532938602777718, -0.0512503498649981, 0.166949517563153, 
    6.78219918445189e-05, -0.0603610659836184, -0.0807099493022573, 
    0.0409336632267886, -0.0327252852908374, 0.128648583220286, 
    -0.0934072059934071, -0.121838333716344, 0.0112013133158855, 
    -0.11562796194475, 0.0245492734759945, -0.16593755760991, 
    -0.00209191163510609, -0.284260934487962, -0.116413606929698, 
    -0.00260485319475462, -0.208541002059431, 0.00298984061270341, 
    0.0652903797620452, 0.0592346354756244, 0.11213341084375, 
    0.182061671252915, 0.136330760570469, 0.104664676567336, 
    0.171712059829973, 0.123317088781821, 0.114657489028948, 
    0.465233052158463, 0.199737950179917, -0.189197907110253, 
    0.0984780814016155, 0.587876654915123, 0.15735377881153, 
    0.0467138152728882, -0.0506212442540825, -0.136771344158846, 
    0.186852481844709, 0.657297631013156, 0.185770428247263, 
    -0.0841305238587368, 0.0605408033784468, 0.636162066214768, 
    0.000795920767353756, 0.0127365319457497, 0.384696212286409, 
    -0.0708869776509179, -0.0836371462925231, -0.0963811817360863, 
    -0.260735778780615, 0.0843962064652615, -0.233669748696493, 
    0.0835173874450983, -0.119700302607912, 0.119696527999151, 
    -0.2186956382109, 0.0553005758891602, -0.10530686436805, 
    0.150846633653131, -0.0544533524692521, 0.0131684042212716, 
    0.0460950730663446, 0.0802372135450582, -0.00193799663310633, 
    0.0631494659748121, 0.0343975852129674, 0.0417833425615617, 
    -0.0724820680228623, 0.0130633444957434, 0.0649327124338597, 
    0.0602979671453404, 0.0873859510863605, 0.117988766711433, 
    0.0912135531073721, 0.103509604680776, 0.12314586929657, 
    0.0296352507939721, -0.00233071222558692, 0.460239258780108, 
    0.200452593048212, -0.0848279966834665, 0.022556086151097, 
    0.331911904182574, 0.516331318759909, 0.319657074580131, 
    0.133065730843639, -0.287686840299224, 0.611598399544313, 
    0.413326442011732, 0.0343743521693018, -0.117876733357649, 
    -0.212737385214444, 0.40214025964373, 0.279902561430452, 
    0.122624585993242, 0.180480720661915, 0.474565033118423, 
    -0.115086329798869, -0.198237293885233, -0.0837341456330061, 
    -0.150179162126639, -0.139525476923656, -0.183293632747316, 
    -0.156852408924909, -0.190273091073297, -0.109820294222191, 
    -0.193830115704644, -0.0985861731252981, -0.0654130231032366, 
    0.066032842627325, -0.00857086706722407, 0.0368187373167629, 
    -0.0937102665315326, -0.0108083666732823, 0.00915690684982495, 
    5.85079734549132e-05, 0.030753351156206, -0.0524150229057477, 
    0.017439366820529, 0.164687861027931, 0.0431936913216465, 
    0.044626101285247, 0.307279509208857, 0.195363963277421, 
    0.0977405612076169, 0.00669807917747652, 0.152928692846368, 
    0.270533676843668, 0.0408970631840737, 0.874608685855069, 
    0.34271000476622, -0.149081581664055, 0.298114478058825, 
    0.77571360441593, 0.142533524650945, 0.129060968230065, 
    0.109077739202231, 0.666980255797612, 0.0553664406533526, 
    0.00258875099901502, 0.0955745392238192, 0.0238751851371518, 
    -0.0391670356458286, 0.054305717057381, 0.0367692643022133, 
    -0.0415100190998562, -0.0503867472517585, 0.13211527463744,
  0.360930000321005, 0.00490525224286693, -0.0784832439205185, 
    -0.0916941067084075, -0.0158147210992065, -0.084693131503476, 
    -0.0923733657668918, -0.0943369348626921, -0.168029951180074, 
    -0.0949862822649327, -0.0513055411605906, -0.0528951908265201, 
    -0.0399377521909643, -0.0562371839827727, -0.0146711907695487, 
    -0.0597174908777068, 0.0212215443098217, -0.0339966752823884, 
    0.0649698828207706, -0.0749837921832716, 0.0230506515247966, 
    0.0647757402097777, 0.0844341863339204, 0.0918380662753556, 
    0.0891093830527329, 0.0820917916710911, 0.0949110162899372, 
    0.158942731294957, 0.132936139379829, -0.147969904409203, 
    0.210891275677751, 0.279159306473196, 0.159797472334337, 
    0.407802229982694, 0.300114182334128, -0.00525549879986415, 
    0.0478499668122373, 0.0350331413600712, 0.799938587340091, 
    0.522318705131149, 0.0273429583255359, 0.000761469769467504, 
    0.149411272366853, -0.101602222203138, 0.306771724032861, 
    0.206295068845019, 0.0451155390605408, 0.36423476355686, 
    0.234275975260747, 0.028252274108137, -0.118580272435265, 
    0.0361092571774497, -0.397727294364964, -0.141745537706478, 
    0.0199652851329006, -0.306923972547976, 0.0841532680917382, 
    -0.0322842082937528, 0.104533759744857, -0.205489934477238, 
    0.0363186234729808, 0.233404916996194, 0.151812705075634, 
    0.131868187427715, 0.260814104314427, 0.276814853049266, 
    0.233279630463014, 0.247488043224341, 0.209270680122969, 
    0.159044276247004, 0.401945411325417, 0.463046142710626, 
    0.231301599989148, 0.0231116136205777, 0.450414256319211, 
    0.594604099410987, 0.208182471543191, -0.108570320880218, 
    0.330762334667625, 0.547367743360415, 0.375620059161934, 
    0.242761648728251, -0.184974181386138, 0.528568017687488, 
    0.417457255672012, 0.0943937161671795, -0.320775323357507, 
    0.185547431837435, 0.485561114499374, 0.0126014646937183, 
    -0.110618103639011, -0.0359770541873951, -0.113039420053863, 
    0.0188484368480784, 0.0693496962853126, 0.422351171562589, 
    0.199819722330873, -0.0433383002212618, -0.000405422548681173, 
    -0.00665059718734776, -0.0842673936940408, 0.05112478331102, 
    0.284403879998674, -0.0777378211965913, 0.202261288558477, 
    -0.100534584063053, 0.146017884427231, -0.0723707612266856, 
    0.172578212061935, -0.213850718946415, 0.107208710884613, 
    0.117233048319576, 0.114529489299179, 0.175961268714909, 
    0.162736349406493, 0.0708572097970931, 0.0825574507719593, 
    0.163735524933674, 0.13684868308774, 0.066530729550614, 
    0.0647076372197275, 0.0258612486077467, 0.0357489297008663, 
    0.0346560757633935, 0.0329568120414973, 0.0497839138010385, 
    0.0226326171115645, 0.0531393215337627, 0.0798396693641477, 
    0.0055705638182352, 0.255208470613303, 0.00562563756491323, 
    0.297002333207799, 0.562155820322306, 0.0298716119227742, 
    -0.134938830084354, 0.28182886312528, 0.220275611845999, 
    -0.0818246059943253, 0.182228044695396, 0.721061117842838, 
    -0.118754126695429, -1.20746655354331e-05, -0.22794316692011, 
    1.18513458483223, 0.526705029422921, -0.116459731938966, 
    -0.0129636018272562, 0.770726904021609, 0.296690163127004, 
    -0.0328952258991378, 0.0655029653294083, 0.179834479402109, 
    0.157420186407939, 0.11746814058718, 0.0590510513080585, 
    0.00333857918275746, 0.0957699509448683, 0.10108083205885, 
    -0.0133344379218455, 0.136106174907392, 0.338367163618949, 
    0.114839855401698, -0.0970318405893891, 0.0190345138298864, 
    0.215090268942395, 0.250701355863558, 0.319723082245774, 
    0.193407591687302, -0.0791832470343058, 0.252339133634353, 
    0.33120998907764, 0.105332921815823, -0.0103494841981224, 
    0.427371038640031, 0.167020790233414, -0.0284293946115148, 
    0.0890587049628345, 0.367872287820273, 0.145195557243634, 
    0.0143210511477985, 0.021181891395428, 0.0412501630790251, 
    0.0455633391523972, 0.0625145183184558, 0.0327766872722771, 
    0.046800447931121, 0.0903873166879787, 0.081584036815133, 
    -0.0490548688099569, -0.00894148402945853, 0.343112311145526, 
    0.140427004959923, -0.0472494190068073, -0.0285570096957826, 
    0.402492822511407, 0.245805365347258, 0.0842794840115902, 
    0.0290012417842805, 0.155611152630648, -0.296226157748248, 
    0.0897115706573121, 0.889105000894256, 0.345422359110071, 
    -0.294371436503285, 0.727829160580157, 0.375046262167719, 
    0.130934346221262, 0.788069109452666, 0.0189774828372631, 
    -0.375828199969575, -0.0797427943462316, -0.12905351701093, 
    -0.15097039748264, -0.125831451258471, -0.0792853633793179, 
    -0.0251782098229169, -0.216452496525215, -0.024351660141151, 
    -0.134785053838177, 0.0943201663691952, -0.0826764284724889, 
    0.0490359672148696, -0.0139436798639395, 0.050218351887478, 
    -0.0526853855400038, 0.0300931179394938, 0.0252192928537866, 
    0.104753422394301, -0.0273824370435991, 0.190633908792543, 
    0.109405020625218, 0.030278718184333, 0.000663505326827338, 
    0.0911781192478514, 0.0939166739851003, 0.356725453132073, 
    0.203276266944921, 0.0138107274461379, 0.127725107547097, 
    -0.0523250019351874, 0.0487545950149422, 0.592445897140597, 
    0.507275045487638, -0.4995400619383, 0.522483668324473, 
    0.716147494208124, 0.525680066660022, 0.980768594637453, 
    0.469390145398087, -0.0671296380114886, -0.127785342059002, 
    0.118773940782095, 0.238300520555567, 0.229942297452356, 
    0.15325126372666, 0.135825436230934, 0.0372603643654891, 
    -0.425285436717132, -0.245259018052577, -0.198056395511925, 
    -0.207479365581767, -0.198701242304254, -0.187822478447644, 
    -0.171677336783511, -0.0341008246100407, -0.156929936013985, 
    0.0629807977156205, -0.268982272659953, 0.0115510674906214, 
    -0.100508044065927, 0.0125990627128061, -0.198701307318217, 
    -0.077012363479328, 0.0368199320929726, -0.142123862851828, 
    0.0326087700794421, -0.110501288888383, -0.086409719117821, 
    0.0108730695288337, -0.0654783076956134, -0.00860019755673341, 
    0.191120917281945, 0.0587243047870852, -0.0207250825833307, 
    -0.0706633536369274, 0.145119025024549, 0.253466219838459, 
    0.0269841536236137, -0.126583310761979, -0.301295991941763, 
    0.976894925177507, 0.0158449564235708, -0.439225387708715, 
    0.178081930027947, 0.575902644544778, -0.101833426305568, 
    -0.210988509620096, 0.0787002540933982, 0.65331158453415, 
    -0.080557479939464, 0.0292275619273745, -0.0408280921426054, 
    0.283615510771562, 0.0995601155789344, 0.215176685996385, 
    0.37983790648846, 0.0205552560066645, 0.367361918434441, 
    0.579491004917612, -0.0461843032099986, -0.081011444392162, 
    -0.11652149227665, -0.06264310190622, -0.159136742384384, 
    0.0289917103657735, -0.0573595526245566, -0.0645627331922178, 
    -0.0865140586770534, -0.0356543635419818, -0.00463200714829914, 
    -0.104568323182085, -0.0125859061705625, -0.0338933006866744, 
    -0.0432704587845461, -0.00829225437047389, -0.0461969524614981, 
    -0.0087425552483833, -0.018532938673293, -0.0483879169615652, 
    0.0515013598700636, 0.0108518406581169, 0.0375915695411373, 
    0.02048817805675, 0.0316337889826202, 0.00533876304433341, 
    0.0136877276370752, 0.0376773435457877, 0.0211234839660909, 
    0.0115449631548346, 0.039962895910944, 0.0200847221160811, 
    0.142714743072299, 0.249586448922774, 0.209461993005111, 
    0.128506416047603, 0.26269647459493, 0.260737816262281, 
    -0.00399199576534766, -0.277805231508168, 0.640324150188581, 
    0.334788919296835, 0.441305246532682, 1.09468310270448, 
    -0.0531482665205269, -0.144548720349205, -0.129245889277614, 
    0.424133556365577, 0.488703888311296, 0.593708374680488,
  0.05179389131563, 0.162000825024038, 0.190940453870053, 0.105046457619574, 
    0.0673816965886995, 0.233932880671857, 0.236087842712467, 
    0.189447068300281, 0.195813859609874, -0.247605023669488, 
    0.553899164437393, 0.3768526994385, -0.112006118271399, 
    -0.0517392023862766, -0.539587807678497, 0.478658387641507, 
    0.430978643949056, 0.0835912952371703, 0.916389246770782, 
    0.376619652520985, -0.207975461755144, -0.0410535103264653, 
    -0.0321945641423778, 0.218598564047836, 0.0710650563102302, 
    0.140814213111408, -0.275398791021535, -0.123868940576756, 
    -0.134770812643549, 0.0884448913551073, -0.345192525738124, 
    0.06591487316207, -0.241684307468587, 0.0921241143448556, 
    -0.243275832514901, 0.0651092671680624, -0.393724884809656, 
    -0.12375069204948, -0.127185223122924, -0.233143250838257, 
    -0.0455897432603865, 0.0158707720037306, 0.0379412757592992, 
    0.066741196085275, 0.0685217680387883, 0.0560743584582867, 
    0.0677167213345491, -0.0923346989281618, 0.215786907397339, 
    0.20188560649605, -0.0497407941224227, 0.238934352877356, 
    0.594692618024715, 0.115195875168885, -0.315396090936498, 
    0.092770555476152, 1.04372067432832, 0.242676885174546, 
    -0.114964923124314, 0.28449662332606, 0.488705630842157, 
    0.0486639026190911, 0.0108197058479225, -0.0387318928420805, 
    0.339535007856875, 0.187258035154692, 0.120593683641315, 
    0.432792645562617, -0.00750132469156115, 0.0300681463194464, 
    0.0392424917454974, -0.215787126382186, 0.164922706711429, 
    -0.160775893913986, 0.162360834318415, -0.279898648761821, 
    0.0768011920915828, -0.357559478843378, -0.0685347185905763, 
    -0.171170615287869, 0.00896560404095681, -0.0280164648573055, 
    0.31066303898258, 0.23560789331084, 0.0721431492108268, 
    -0.0362464182051175, 0.221541532437235, 0.390482081308575, 
    0.281305611923419, 0.204285937631724, 0.258614793518723, 
    0.273042818186044, 0.253884519023754, 0.39002449996677, 
    0.529614069575257, 0.378825025683, 0.177432583058506, 0.234057179122499, 
    0.551181223511935, 0.391314166632319, 0.123495036494495, 
    0.0750749662176148, 0.472392442246515, 0.434377084647579, 
    0.0958690309874953, -0.198060387430494, 0.0835568082875306, 
    0.507515887000834, 0.0897688806491099, 0.0388732050974665, 
    -0.163854596958953, -0.136869478656069, 0.413838550160042, 
    0.381547778696628, 0.119913230331203, -0.00515041258765303, 
    0.00592975866299124, -0.273743922683359, 0.545418946441904, 
    0.187415922248662, -0.0859048705895053, -0.0731094094486037, 
    0.0883803416009408, -0.112854267428342, -0.319971027312639, 
    -0.172822177650778, -0.149768076008971, -0.0805343206706701, 
    -0.0930429999298953, -0.0888206563704253, -0.0890258505610052, 
    -0.100845449709956, 0.183133984138072, -0.110088459836915, 
    0.179513541054967, -0.332179735235598, 0.0683346958493179, 
    -0.294943846103725, -0.0289599219891378, -0.304914386150103, 
    -0.131997841976705, 0.0543349864219303, 0.122511260175401, 
    0.0649457758189056, 0.13300201438277, 0.235469887268378, 
    0.188249945344513, 0.113630692399885, 0.0814303767324431, 
    0.116448876232752, 0.242397512681921, 0.275863139800689, 
    0.252362809555582, 0.243460846348876, 0.254628709225056, 
    0.234898054980568, 0.187801740912175, 0.17842298028409, 
    0.258050498810784, 0.289141242015291, 0.213901912732598, 
    0.15947046081637, 0.132215160965267, 0.138196015935195, 
    0.170656531454356, 0.151857895566864, 0.133184526687026, 
    0.191286964831759, 0.112807052558062, 0.282054719491351, 
    0.312664932578934, -0.0139620204764102, -0.140971242619658, 
    0.0681851653739083, 0.480354139064436, 0.505393762785504, 
    0.518209129378338, 0.230320646359403, -0.11071231404768, 
    -0.262844875229039, 0.470935237641055, 0.483646268687631, 
    0.178179101546858, -0.234721124668835, 0.196339798195107, 
    0.165349346952933, 0.190433066253654, 0.549841715076817, 
    0.247328016429009, 0.0399062750254264, -0.0423058682758864, 
    -0.182008888351169, 0.0834319892852427, -0.0873366673986419, 
    0.0285853977423651, -0.0961420011044172, 0.00484387952397256, 
    -0.179253621957992, -0.0869706447511526, 0.160121189898718, 
    -0.135007035392206, 0.10519520368568, 0.42498028755975, 
    0.0391254001922355, -0.0510479377288701, -0.200050941344217, 
    0.211833636971835, 0.466564064077901, 0.332048993840093, 
    0.158018521795905, 0.0382773492664656, -0.0257197759125036, 
    0.546781463827316, 0.28745525334386, -0.233605122822085, 
    0.206468864010735, 0.924473897553527, 0.169133087474038, 
    -0.163896795475822, 0.136239773576153, 0.640135025622966, 
    0.197745952075525, 0.0387898437204733, -0.144268744929889, 
    0.150868888025105, 0.520923709446052, 0.123243552304899, 
    -0.0163101130180286, -0.169193032120321, 0.15015335691816, 
    0.479352219901081, 0.0677796244295656, 0.0463999837922586, 
    -0.316948215132016, 0.50329173836039, 0.234909547180133, 
    0.0192354491999494, 0.459183247933221, 0.0725651194573968, 
    -0.114993878517914, -0.210389344202059, -0.115178082940717, 
    -0.0198572136808577, -0.198691994331557, -0.0252838705676628, 
    -0.112484848743406, -0.0639084951119923, -0.102915475038519, 
    -0.115591523637231, 0.0491372829361644, -0.206620737210832, 
    -0.0179843408278427, 0.000394930341667862, 0.167256586962644, 
    -0.154788458145294, 0.0983108585817194, -0.264312547471198, 
    -0.122459909214737, -0.0571427501259451, -0.343181013548446, 
    -0.0737765926058369, 0.0318389166527641, 0.0238046911057674, 
    0.0393261688711123, 0.133379972096734, 0.09864873699631, 
    0.035310721997929, 0.120639937451062, 0.18589210311679, 
    0.0550899812097286, -0.0792634946668584, -0.0165273497604827, 
    0.493872267515197, 0.221857983995752, -0.0200799673064579, 
    0.333934699512944, 0.323643609971778, 0.159381371854182, 
    0.62572332718349, 0.399506750736729, 0.0200668624882237, 
    0.00169866157363496, 0.0927725110095444, 0.562347508856909, 
    0.589374241714612, 0.142637137319876, 0.206230261125221, 
    1.05329582434487, 0.105397180373993, -0.066179352744485, 
    -0.224673468890964, -0.164623342196671, -0.118144020453294, 
    -0.195507725974261, -0.119323404190881, -0.212184509640924, 
    -0.122943208444429, -0.162453178572099, -0.129922416466924, 
    -0.130937053622246, -0.105995745711962, -0.0107810688881469, 
    -0.0238636830497165, 0.00146189146531657, -0.129931665528522, 
    -0.00456278409005261, -0.182631817051931, -0.120683264221861, 
    0.0347659866260368, -0.0992762863180097, -0.0388447175720964, 
    0.0457517078640039, 0.0648690337528399, 0.0858357648060804, 
    0.0863460008847116, 0.0555862826160457, 0.0582410122264042, 
    0.131272883728725, 0.0756755254808672, 0.0222898314737216, 
    -0.103644243196557, 0.323079218676176, 0.283300066557296, 
    0.0807906719230919, 0.00181682363739137, 0.0304820710333102, 
    0.224600831630339, 0.714836110296294, 0.260803198999457, 
    -0.24159822974544, 0.415047543585539, 0.418550928157117, 
    -0.16575928292647, 0.301432483171627, 0.625360766911374, 
    -0.156865516796402, -0.365867653777249, 0.205682177839071, 
    0.281200231105066, -0.0596323151728956, -0.241249202807126, 
    0.104079909890222, -0.161528249065627, 0.0916874713252935, 
    -0.217746639145864, 0.0588095412005578, -0.24749127291042, 
    -0.0325956738940865, -0.207321235134561, -0.137540090230758, 
    -0.00426601542853043, 0.093788436304838, 0.120309169992474, 
    0.0921434273693409, 0.0248375357780793, 0.0445885377535811, 
    0.0657404820903583, 0.127112334793672, 0.133130925678086, 
    0.0463985201393063,
  0.445402847405252, 0.156703870034046, 0.0657219497790163, 
    0.0860726264459704, 0.0892624591093214, 0.231693856283294, 
    -0.0659911748134035, -0.0816930942755171, 0.0114373859649932, 
    0.187657908241419, -0.102932423177633, -0.0352111804264537, 
    -0.181496948709365, -0.0214197821221536, -0.0827483426822756, 
    0.0504961938108375, -0.277794951217133, 0.0527031135894952, 
    -0.353750042019011, -0.185132562371176, -0.0214280713179985, 
    0.0532122468557781, 0.100400301006321, 0.157723979798481, 
    0.191911749185329, 0.150297044750699, 0.159095038441517, 
    0.281588800070447, 0.20717737505867, 0.057213971230776, 
    -0.108565326362787, 0.36974702501269, 0.572168124142867, 
    0.115972606568587, -0.210195581517783, 0.063327360875359, 
    0.726751494811403, 0.00166639093922227, -0.172690163756361, 
    -0.0635783446445174, 0.546335869813909, 0.317187933677531, 
    0.215325129229748, -0.275581203289004, 0.355790991410888, 
    0.382688787621669, -0.0956182830753915, 0.245065382043494, 
    0.811242671739539, 0.18974306155419, -0.101501205304398, 
    0.225672123966838, 0.188263132785744, 0.177884233512186, 
    0.575257762328583, 0.285706877028773, 0.0861004291067342, 
    -0.198420716762747, 0.269695158175666, 0.317045492158243, 
    0.0959246425221346, 0.167580463660558, 0.13141012476484, 
    -0.129670120062049, -0.0278664659370931, -0.0534683468641565, 
    0.148799339599315, -0.00192168584672378, -0.0325750413580884, 
    -0.00210974654755794, -0.1183290429797, 0.0507218449626579, 
    -0.106682738414613, 0.00839173887886767, 0.0192638891569602, 
    0.0726878055225142, -0.101007663580568, 0.0409225888249634, 
    -0.0782405763367219, -0.162593010698689, 0.210983943365522, 
    0.09206406232737, 0.0248678464817492, 0.0856099328961956, 
    0.249213966684612, 0.13095468377472, 0.63792622030963, 0.251402438949339, 
    -0.267734548566736, -0.271747266837992, 0.130706821584067, 
    0.657367602669584, -0.349133006872214, 0.178616528391784, 
    1.08719988227258, -0.0927935930715949, -0.386841567414859, 
    0.0552270966684414, 0.777582490205858, 0.152068366700616, 
    -0.0666921573226914, -0.162545094215085, -0.114472201097794, 
    0.450485643787631, 0.324711090316866, 0.0399087840281924, 
    -0.0583694197830828, 0.00896179665671157, -0.0883798662987695, 
    0.184498124582986, 0.425728031505643, 0.144264353864306, 
    0.00952498881939767, 0.0784310152730506, -0.211925881637342, 
    0.311740256072272, 0.20364890883952, 0.0732168609599703, 
    0.0666162510213901, -0.200806037457753, 0.0023997426430979, 
    0.366968718029689, 0.296733722331393, 0.110754359658581, 
    -0.136947291983634, 0.0328836704865867, 0.384536435264392, 
    0.2280196851655, 0.104191926724141, 0.0648640140614144, 
    0.038314158751447, 0.141407008471407, 0.328972644633697, 
    0.258573270560359, 0.109200180609595, -0.00782722660355457, 
    0.290162154143567, 0.299811573191241, -0.161082017313015, 
    -0.0896150470529593, -0.110035373899034, -0.119548763338625, 
    -0.0361613601800024, -0.153483062308265, -0.0437491211334848, 
    -0.140914813246527, -0.100444618191597, -0.0540585767365375, 
    -0.113919027907096, -0.0566700396163163, -0.00440167828495415, 
    0.0296622323885612, -0.0402295787427889, -0.0061050919622291, 
    0.0192419081647222, 0.0288280078458173, -0.0332544766458457, 
    0.0124939758294356, -0.0573267637751603, -0.048690674157114, 
    0.0252688945263978, 0.0841056214418832, 0.0578156590903864, 
    0.0622114617530826, 0.132400213901699, 0.0953841970860303, 
    -0.00260145802384174, 0.23139220265587, 0.120085891395064, 
    0.168877292661809, 0.552322634475711, -0.201403185778309, 
    0.587575281465747, 0.529882087674523, 0.0748363615806496, 
    0.0129883099238301, 0.60403672369089, 0.356105906636329, 
    0.392128145068036, 0.717613868832661, 0.161703430640462, 
    -0.0103561150380475, -0.0293406827779733, -0.00171225834206598, 
    -0.0578556835360152, -0.00454789299266425, -0.190933917380788, 
    0.0556814274793942, -0.22811318783756, -0.15038135676095, 
    0.0376445802738913, -0.340708392696278, 0.0491390317088795, 
    -0.193199767778164, -0.110004733290432, -0.0335536408158988, 
    -0.00833532802207487, -0.201505791545716, 0.0649584808447106, 
    -0.308022032328489, -0.121309994516012, 0.0384284102944578, 
    0.0666922189006737, 0.117390606441681, 0.156957651762471, 
    0.119610777669656, 0.0946408876048426, 0.102941384725288, 
    0.0999807265858684, 0.0838264045362535, 0.178214675351428, 
    0.215648539231557, 0.225994213122699, 0.242656506709389, 
    0.222778693657158, 0.177501893204609, 0.244350159699469, 
    0.337301046986678, 0.187366758538159, -0.0630622581483769, 
    0.432075119266262, 0.365217780783908, 0.0323293650976762, 
    0.123531215468879, 0.643323275270814, 0.287964533384587, 
    -0.12770236669032, 0.679608333712393, 0.351885563929201, 
    -0.0878803262275683, 0.567088239212136, 0.468922989899757, 
    0.0635194320341428, -0.32295737106424, 0.466741035314937, 
    0.693624442974025, 0.332944649758434, 0.0692932427512113, 
    0.797772430289551, 0.300076732206936, -0.091116591604832, 
    -0.217120517183553, 0.0579175567573943, 0.0782907937011623, 
    -0.0693283335573844, -0.110922828966936, -0.074294085964321, 
    0.0079339760786708, 0.0460864523055103, 0.162902711984261, 
    0.0812969013224179, -0.0200342901456442, -0.0514710387824481, 
    -0.062276880538177, -0.033132104062313, -0.0954169712293668, 
    -0.0303613536181755, -0.0912999341427085, 0.0248985784480371, 
    -0.114519654216431, 0.0239992479488815, 0.11161964393604, 
    0.0937894952267083, 0.0730548436616306, 0.147763866343733, 
    0.189292716303477, 0.137066104353656, 0.099348125520846, 
    0.126500673031808, 0.175173110328331, 0.177011327637749, 
    0.131541378012972, 0.0947200196578417, 0.113780118328357, 
    0.0908941956551095, 0.0711691538291573, 0.0870910507653201, 
    0.129410648498141, 0.124494202758535, 0.0365258321754999, 
    0.0872492074229633, 0.255079717231723, 0.187130983700668, 
    0.0402231419355468, 0.0326947741266881, 0.394171757210302, 
    0.246262780305819, 0.118805162945012, -0.236125775307138, 
    0.456111102174905, 0.359230398228041, -0.110373445972855, 
    0.377681151560826, 0.483560479646397, -0.0144630097927691, 
    0.386241989580075, 0.611070987903007, 0.130435365994114, 
    0.0952966547863061, 0.396175205257836, -0.0250096788633598, 
    -0.0547352937412098, -0.177500829107243, -0.0601355626796626, 
    0.159545832412809, 0.0844443165836237, -0.123458630932899, 
    -0.116168232615122, -0.0695802494443913, -0.0396880592260271, 
    -0.126772163936861, -0.420690980289973, -0.0550966407920234, 
    -0.00730952775565541, 0.129276432133206, -0.249154827399455, 
    0.151723577896015, -0.17971354687942, 0.0348680596284517, 
    -0.504937816695017, -0.0950494855580044, 0.0250514367546665, 
    0.0262616548009812, 0.0640109978124783, 0.108544384194177, 
    0.100186779930598, 0.132088248603016, 0.171465177623191, 
    0.0985725654864468, -0.156576893561272, 0.31507135246755, 
    0.448313182437535, 0.132891781241059, -0.271537429719623, 
    0.196467096512643, 0.609403219858495, 0.046068839730957, 
    -0.12242123709913, -0.0304490877068365, 0.633319866375197, 
    0.0182988720567603, -0.108143792042238, -0.0848629391770434, 
    0.586577138124272, 0.221223049869834, 0.0869671472688185, 
    -0.0296082528377681, -0.142667216119179, 0.649198512303828, 
    0.131301357818275, -0.0573167931664016, -0.045310572540942, 
    0.470018107677362, 0.0811154214060044, -0.111782065273571, 
    -0.192276468005693, 0.499199606956571, 0.466162399854014, 
    0.224423537201606, -0.0429075227402928,
  0.458500421788385, 0.459541216997255, 0.374842135634717, 0.330443704265065, 
    0.265906837327605, -0.412130384527005, 0.69805697545425, 
    1.11629352570972, -0.407764416449646, -0.203634169261666, 
    -0.192858624892072, -0.303722264535698, -0.165986670850342, 
    -0.0604209239535829, -0.102828256551357, 0.336614620236183, 
    -0.283142185480601, 0.166152320125282, -0.30209521850502, 
    0.00809414695507155, -0.0837359976136862, 0.10535590442589, 
    0.137996789477156, 0.17177655827938, -0.037998062545294, 
    0.141604932683536, 0.0604826857619764, 0.14400820062915, 
    -0.0159000092433837, -0.205224964267114, 0.0108710633283827, 
    -0.137502768233636, -0.0961732036783432, -0.0992650993304225, 
    -0.0900033890547154, -0.0808479919984661, -0.0801649328715152, 
    -0.0619757038753807, -0.0876091529014889, 0.191308628835264, 
    0.442095776578637, -0.0738136219464198, -0.29133013609763, 
    0.149170828816536, 0.303530666591032, 0.666328155754867, 
    0.647226683182172, 0.183635098287277, 0.0647795032637377, 
    -0.407381865947198, 0.11984335475008, 0.491896523286706, 
    0.214071763921797, 0.0591066860186533, 0.0654628428095919, 
    -0.318191205489165, 0.438931985961982, 0.389789302726459, 
    0.159492417642281, 0.364763954295763, 0.336219084261999, 0.1401785072644, 
    0.0505615208891137, 0.0187558988777865, 0.00519256235143537, 
    0.138747632567724, 0.152087954936379, 0.0552876719357533, 
    -0.0180816174041373, 0.0810093567465783, 0.407217929613148, 
    -0.044734697985188, 0.173102887878334, 0.597752155551575, 
    0.19284424970351, -0.0966766630216474, 0.429041269441858, 
    0.443727244328833, 0.221624837587464, 0.139382662128148, 
    0.167095579231328, 0.181528284981437, 0.10518156701926, 
    0.095530671727938, 0.0978653517268, 0.0361188905890088, 
    -0.05111030446009, 0.107469933711978, 0.106612739983538, 
    -0.0242363715290295, -0.0646282554454402, -0.139061343929854, 
    0.0174209308415944, -0.0552636288225632, 0.0294646254129694, 
    -0.0926180282040521, 0.0398917100354079, -0.0971508084207113, 
    0.0160497883072104, -0.182927816085746, -0.0292710809556011, 
    0.0233420266225695, 0.10293983470895, 0.0909438491565469, 
    0.054487298474165, 0.0584346905427354, 0.0179505334722849, 
    0.362686192855432, -0.0139919132974326, -0.131527940711889, 
    0.111671813572176, -0.0235364143187394, -0.042783611799977, 
    0.95432147949481, 0.233609338250399, -0.30736746876609, 
    0.0858090068674295, 0.855997230675418, 0.36583301745896, 
    0.148937987665215, 0.380756329065077, 0.302255265499063, 
    0.0871212289674897, 0.0904580277830391, 0.216057432629474, 
    0.0367744393137584, 0.377236652497403, 0.00341258362465127, 
    -0.0943056006596823, 0.099899885028199, 0.243549876908574, 
    0.169428658695823, -0.0928500007722987, 0.252037350130133, 
    -0.255528394304238, 0.0774779589840211, -0.170760598090804, 
    -0.011791847185094, -0.459370899104603, -0.157946047312835, 
    -0.040862964354295, 0.106098359646571, 0.0497979982388603, 
    0.0504494093338494, 0.107862681009622, 0.0788162705022761, 
    0.044420902273944, 0.0870813916514728, -0.0157146214248413, 
    -0.0256082049601767, 0.115518212340617, 0.0983613489892824, 
    0.0693076268946475, 0.156626413816611, 0.203015917964224, 
    0.222164865406886, 0.280523939490351, 0.107371830078405, 
    -0.086280249661582, -0.150211928348023, 0.508136887874375, 
    0.302096564276547, 0.12066843641018, -0.265718494716079, 
    -0.00275793739695175, 0.606217433707017, 0.100550484822736, 
    -0.0459680035409758, -0.115518620712016, 0.473010928684346, 
    0.254790376097043, 0.0516783943405797, -0.0590549228968377, 
    0.103065924446246, -0.142716047053939, 0.354368804033402, 
    0.236946634891283, 0.160111415901415, 0.365843154749534, 
    -0.103125182786705, -0.314986597770943, -0.0528094326487933, 
    -0.189992939916848, -0.139953627851817, -0.150348523224184, 
    -0.167610988191116, -0.133672945067651, -0.128855163182282, 
    -0.108672161236131, -0.139720730194744, -0.00268432378692141, 
    0.0335594145751389, -0.0991057279232241, 0.0146806108990945, 
    0.00352074770801131, -0.0561218281325958, 0.0787139252844742, 
    -0.0178479280535622, 0.0300169184475601, -0.0451330782392963, 
    -0.0273146399728053, 0.106416592729116, 0.14440707981802, 
    0.0719031410176198, -0.0210589782716277, 0.138454299773927, 
    0.298492999942098, 0.0426468838619422, 0.0625941393569798, 
    -0.312301218161875, 0.17230248959662, 0.397791212788465, 
    0.471187282878715, 0.323145329574831, -0.0018071178518488, 
    0.685391914887218, 0.206843348718894, 0.0526285527313647, 
    0.101835779638007, 0.623954565056922, 0.0367811725412759, 
    -0.00932020446009924, 0.00494396061950543, 0.124169397623044, 
    0.135281308666795, -0.150826046688077, -0.217301695350103, 
    0.0036258105719589, 0.0130520314973453, 0.20330291015196, 
    -0.173360963770144, 0.202549788322427, -0.178577206819378, 
    0.100260500536971, -0.0656234039513158, 0.0851003859317901, 
    -0.402465211748535, -0.0443664999679257, -0.173483831312284, 
    -0.252854422352593, -0.0056615918971263, 0.0503421664713961, 
    -0.00308085023600585, 0.0342278136569328, 0.0600642845441072, 
    0.00949182062716458, 0.0396164652777384, 0.0623909243772398, 
    0.0568047557436727, -0.00256042920290023, 0.0813243976357157, 
    0.113952457266454, 0.129402458836033, 0.178692822877661, 
    0.167566567638041, 0.0772318565098982, 0.166398516210669, 
    0.39336840905476, 0.0997350733696297, -0.164708547455658, 
    -0.0297613179916842, 0.480548575577534, 0.262721152325703, 
    0.0843121947198545, 0.0414286194873045, -0.229676181486262, 
    0.491155132543779, 0.355985206455894, 0.0939987206205276, 
    -0.00078984373280494, -0.124112706661021, -0.0227741816530554, 
    0.538498426068385, 0.226697642284893, -0.0191519812751011, 
    0.0861348217769003, 0.287179571438929, 0.419012246125237, 
    0.0337968477400964, -0.125684641630437, -0.306892312777579, 
    0.148509918246252, -0.31251812772107, 0.0829167982482933, 
    -0.328957843910461, 0.0310750122520399, -0.332757342476451, 
    -0.0526135128124756, -0.238353902079881, -0.123626105101186, 
    -0.0440856000358472, -0.00242028058131043, 0.029202412314662, 
    0.0582996655528902, -0.0132990476092152, 0.06761161646995, 
    -0.136095450475341, -0.00253440398779674, -0.0280200964097338, 
    0.0150753230314229, -0.0468303484560635, 0.029985405267733, 
    0.0738783486225941, 0.0261265670526126, 0.115966398602122, 
    0.106760681497975, -0.0236480711587179, 0.302926428659957, 
    0.246118982580781, -0.372768993502369, 0.194354335993638, 
    0.603372540139715, 0.00477240037096484, 0.220216645529317, 
    -0.0608809755183607, 0.746821689134516, 0.310086139566383, 
    0.243638194688206, -0.022935079760856, 0.656700060751522, 
    0.240308956575706, 0.1057910071611, 0.152923000840077, 0.167835850949319, 
    -0.0704423621495121, 0.119831825378983, 0.290905430193955, 
    0.1573388718545, -0.154171244919632, -0.243100088247241, 
    -0.29647732467855, -0.132092472413969, -0.155344667938481, 
    -0.262439662708187, -0.0456265317326796, -0.242944347529587, 
    -0.0437110441528546, -0.191714905559193, 0.0591134531488408, 
    -0.222576124870904, 0.0744576259139774, 0.0169711132064797, 
    0.0453303486565684, 0.0378679183180246, 0.0467120166954568, 
    0.00865252276888273, 0.0391629468310996, 0.0183913411382739, 
    0.0186771691440262, 0.0305570135256475, 0.116370263957659, 
    0.013886282621243, 0.22679777303548, 0.264959373755699, 
    0.120273638252957, 0.0051454666977999, 0.250575222738176, 
    0.254540528979719, 0.0422808795033005, -0.0394885110972731,
  0.0639759419322223, 0.0316224652193412, 0.0584993605614361, 
    0.053152213157828, 0.0572118907105225, 0.0346504790665971, 
    0.0410285805246133, 0.104573271695789, 0.0700185994604933, 
    0.11421928660257, 0.390037271491711, -0.0150306542538616, 
    0.317244334231071, 0.322122005527068, 1.010516015161, 0.589670406456476, 
    -0.0881966079315624, 0.603726303895552, 0.440951252968132, 
    -0.197214463291767, -0.178192647549013, -0.0384226135780141, 
    -0.160782539195647, -0.0864137624665745, -0.155725036774801, 
    -0.0910715242211957, -0.119004668960483, -0.100369082831119, 
    -0.061829764014824, -0.0845533934742244, 0.0739037912582046, 
    -0.0435571906632717, 0.0691277677982136, -0.0462229939385315, 
    0.0416076429815703, -0.100325386605503, -0.00575949838537375, 
    0.0172619717966305, 0.0567350817825273, -0.166918143743418, 
    0.0362134664902147, -0.133801173598101, -0.075236048662898, 
    -0.0826229054214065, -0.075669208291354, -0.0963153317339354, 
    -0.0675897130461434, -0.0924204474362139, -0.0456148743294068, 
    -0.178321250400186, 0.0828004703593435, 0.326078168485233, 
    0.242399710835096, 0.199788941831434, 0.776078271075446, 
    0.320667859352304, 0.102849508987366, 0.264960885489083, 
    0.213546567384783, -0.354550276159839, 0.270523284776615, 
    0.302006839541135, 0.334275414792168, 0.604873059393032, 
    0.148320003265536, -0.0600815141819913, 0.212385234625137, 
    -0.35181588003263, 0.798654961753761, 0.273864781351818, 
    -0.289623441252492, -0.207493214682324, -0.13546780296113, 
    -0.106280122577316, -0.142248369092959, -0.0529058847813206, 
    -0.0915481989365103, -0.0745168987094683, 0.00952781962337818, 
    -0.237828394736401, -0.0932679962781843, 0.187177546018089, 
    0.156023904168305, 0.0651886628613286, 0.160288761485789, 
    0.239697303243523, 0.155856725869709, 0.0831276769517217, 
    0.160299149288995, 0.222007873619161, 0.181012401551405, 
    0.144010374121788, 0.144362886615075, 0.153712194089261, 
    0.149425823786469, 0.135029382800443, 0.166974752954436, 
    0.221429732143925, 0.158120241478253, -0.0842565094155107, 
    0.350549402553533, 0.294607787160305, 0.103314382147601, 
    0.329862879139161, 0.323594135262915, -0.0624004683299697, 
    0.116481946101988, 0.483238143008124, 0.455931463261918, 
    0.390655555419176, 0.534586824272503, 0.40587750892046, 
    0.0368400967142599, 0.617048258568421, 0.137101953426298, 
    0.0302083252362864, -0.351458304681725, 0.0022593894256277, 
    0.698781051438357, 0.0863750338377846, -0.127708069113563, 
    0.0509652681790848, -0.538196569095004, -0.109709947247749, 
    -0.147056394899064, -0.296284136442714, 0.0632476072356408, 
    -0.336679807254743, -0.0170779014915713, -0.212416171808112, 
    -0.0727162760751197, 0.0512133045362612, 0.195707751696454, 
    0.175841163244132, 0.0922359758313761, 0.123147748934147, 
    0.102758398656967, 0.118257608464187, 0.098780774748506, 
    0.0543913493423005, 0.130245881119231, 0.219410981538761, 
    0.205414440885685, 0.163266215747893, 0.176408288722881, 
    0.01111208931911, 0.251260151582498, 0.480140830500089, 
    0.169882849960917, -0.148215401682475, 0.472869577512146, 
    0.45131065223428, 0.00767808110988974, 0.393221470482384, 
    0.421432733102061, 0.253180963863876, 0.686446572976433, 
    0.548431564844807, 0.135972286690786, 0.0742624309441587, 
    -0.246859861711826, 0.193048385955993, 0.335497548849962, 
    0.158617201663765, 0.0723750701352758, 0.045178309109092, 
    0.0347206488398254, 0.0401058303333879, 0.0462920455798313, 
    0.0226415953911667, 0.0821908444665085, 0.10824031136071, 
    0.108892399495785, 0.130002927011671, 0.158942268282398, 
    0.122144532879199, 0.0708363963757259, 0.115719278842532, 
    0.131470169012059, 0.0696950151903777, 0.230185986797531, 
    0.432254190691592, 0.288112433839843, -0.0891579830260278, 
    0.282251220775622, 0.124999766224714, 0.536896394417531, 
    0.86123608928256, 0.139985393990844, 0.110986245936095, 
    -0.320946628875725, 0.548578440110035, 0.220691689502313, 
    0.187288749218168, 1.14498121976223, 0.464344571296273, 
    0.114121196048925, 0.0465475008238711, -0.435690670623314, 
    -0.362288554226386, 0.545118653175753, 0.458121014515417, 
    0.0420858464803884, -0.205481326077859, -0.0211432882649671, 
    0.396854174053814, 0.213108167728415, 0.103198927073032, 
    0.156349236719234, 0.179943388464272, -0.0524150399173096, 
    0.349753643675633, 0.683753645621152, 0.0762392003855381, 
    -0.0720877611689375, -0.118400810645292, 0.301430087700201, 
    0.341003525796233, 0.161254604650641, -0.189240404577525, 
    0.269419108337464, 0.442746487011322, 0.107846802041083, 
    0.133757654448241, 0.180858678376746, 0.0478397452293578, 
    -0.229692731494012, 0.49990457399742, 0.142005520457051, 
    0.0343447119337768, -0.0654005683313153, -0.137549653767408, 
    0.0469404148961984, -0.101828146440915, 0.0358394212468894, 
    -0.220033680661794, -0.00553789875217039, -0.117551756924965, 
    -0.00583185832693706, -0.203335984936552, -0.0381220083979965, 
    0.0841562452861227, 0.155666103833417, 0.10636880242313, 
    0.124597957852621, 0.289530548259978, 0.31701855986898, 
    0.213496247885833, 0.120808169939314, 0.0900489463298507, 
    0.27569340696899, 0.320292465416409, 0.213977382055979, 
    0.274102062527837, 0.480577143779712, 0.337142196317017, 
    0.117989102037552, 0.0921765054300606, 0.457429097458852, 
    0.423382293192103, 0.220563661518585, 0.128413030665152, 
    -0.157809279362734, 0.518475528583553, 0.317499767968382, 
    0.100148266447673, -0.0776753242707865, 0.293822188480684, 
    0.309332152960151, 0.103357692133169, 0.469192898384537, 
    0.569890685002414, 0.236087069948934, -0.0135705432558815, 
    0.890464549628938, 0.0644653077828405, -0.152551374295503, 
    0.184441282973404, 0.554141616331285, -0.0779218636548805, 
    -0.109691708239522, -0.0468244317464067, -0.0995261309376218, 
    -0.0678314632592179, -0.0683611078697603, -0.080069856779918, 
    -0.0273205711547668, -0.0658162211832751, 0.0487895990966286, 
    -0.107624285538583, 0.132992405171764, 0.100343831790647, 
    -0.0312797595676675, 0.163707373462487, 0.382721367713681, 
    0.169529305052771, -0.0693317967084177, 0.422701366903371, 
    0.357871104912684, -0.452722141352199, 0.40212540800829, 
    0.732405435944025, 0.320362124134905, 0.146881953919464, 
    0.117016118331957, 0.211751087647908, -0.481831200876413, 
    0.373747604797125, 0.73057994293445, 0.610806606075878, 0.5082060022891, 
    0.113545191989197, -0.158799370599212, 0.0610781999114857, 
    -0.187267552979942, -0.064747630143399, 0.239942936561068, 
    -0.0141283580461712, -0.098515075223624, 0.115177711368027, 
    -0.133606368249124, 0.121647192450724, -0.373465567375159, 
    -0.163721741593783, 0.00183558693105405, -0.207607739367562, 
    0.0348504183495728, -0.217065291088915, 0.00597334988750092, 
    -0.115107902659557, 0.195955654112519, -0.100272012277799, 
    0.0104943572256569, 0.490101302423436, 0.14278819609363, 
    0.0196348688475178, -0.124877780051659, 0.293350261566621, 
    0.319944470903629, 0.148033814547548, 0.0916598863064143, 
    0.282250595206362, 0.388040609309034, 0.353699079968593, 
    0.34289076141192, 0.302454807182506, 0.18255969760636, 0.15097241191748, 
    0.394400458523972, 0.298785648556293, 0.0502624034064985, 
    0.0301825381477042, 0.0378297661941928, 0.0200227370062459, 
    0.025559702505682, 0.0204972930282452, 0.0218308435259246, 
    0.0312236374429112, 0.0249787571461632, 0.0168734214166693,
  0.237447284680969, 0.0256774555683525, 0.00147523671220097, 
    -0.0464159390736053, 0.112010086647447, 0.0132510467759807, 
    -0.00400555787090488, 0.207729566493197, -0.0107689529126431, 
    -0.0503000030920472, -0.0165193318586489, -0.145641071366694, 
    0.0646993176581607, -0.0724331318912238, 0.0517649522920689, 
    -0.162426965022524, 0.0315454077957498, -0.120961553694872, 
    -0.00342451424461354, -0.175999718785348, -0.0607180177364188, 
    0.0245136133990986, 0.00856670979977448, 0.000365733064744661, 
    -0.0547431635309086, -0.00123987772789462, 0.0221834642398381, 
    0.175065728289832, 0.353604356002505, -0.163715501491922, 
    0.607843835040769, 0.319927130105113, 0.0226203557937055, 
    -0.0452651154197981, -0.310144395980083, 0.586456887784871, 
    0.416310065508589, 0.139977124459406, 0.565915391125939, 
    0.465288502020599, -0.23909421395139, -0.206966922669884, 
    0.663405786845687, 0.624389433330602, 0.373998122077541, 
    -0.0345586123710474, 0.698523623490378, 0.241244860966184, 
    -0.0715352435584157, 0.10897423684685, 0.500604234257176, 
    0.241753114357794, 0.0604597058373664, -0.104267530500835, 
    0.000774622327419414, 0.379451396767067, 0.0763319629155219, 
    -0.182261854636928, 0.0214832071105001, 0.615806201045162, 
    0.118132963102886, 0.0781746378582033, -0.346773691033969, 
    0.642652782290084, 0.225620948910712, -0.0888502421861796, 
    0.00366767861033669, 0.179532054109241, 0.613474257398777, 
    0.691414794985303, 0.273175913018385, 0.104294915421124, 
    0.0652249235791366, 0.00700331823845309, -0.0573043618631437, 
    -0.0468246664573617, -0.0173682764854722, -0.109941019307014, 
    -0.0574646712507842, 0.116581905131031, -0.0310293614521409, 
    0.0679833937505782, -0.0528024197553428, 0.0611805482403023, 
    -0.0950259381892691, 0.012089923109542, -0.123740836680054, 
    -0.0453992785918942, 0.0967394202967916, -0.233601831421548, 
    0.020112676111174, 0.320710594103676, 0.0505694292236611, 
    -0.0635189846694679, 0.144494292674068, 0.257444937205535, 
    0.44842869817631, 0.364669127376951, 0.0623110311637534, 
    -0.073153375420968, 0.0812327012264315, 0.226316911600865, 
    -0.214983878376008, 0.329899496835123, 0.710662460270583, 
    0.12878501574227, -0.155737976779357, 0.335304922208777, 
    0.277730840382878, -0.0116709632169901, -0.0977178680261029, 
    -0.176903472074397, 0.0531374689873029, -0.102591371585429, 
    0.0353860497167385, -0.152684912934859, 0.0233751696395159, 
    -0.10711130270329, 0.0250373262250906, -0.184921923906293, 
    -0.02136528443273, 0.12100566764243, 0.0617331596280341, 
    0.0233251508663036, 0.170411598833478, 0.348606205433106, 
    0.137880477328289, -0.157184631035882, 0.115063556883262, 
    0.352551771422649, 0.124282786205772, -0.215154903707806, 
    -0.163755775253093, 0.696683793129195, 0.464859642063657, 
    0.307645401082348, 0.30103172466501, 0.124112421731056, 
    -0.342838042202618, 0.449816895607312, 0.359231566002271, 
    0.264625591905841, 0.476943347056942, 0.294443022000422, 
    0.0759180799992915, 0.102940335941836, 0.316453750300079, 
    -0.0100838796585355, -0.167680459724151, -0.0475091551136197, 
    -0.223310333903688, -0.258283201587218, 0.09919166773154, 
    -0.0912562838493788, 0.11727879623072, -0.208115567219092, 
    0.0207090250694716, -0.178160105426913, -0.0202632697499407, 
    -0.270732495093063, -0.134153128153539, 0.13718133953737, 
    0.012563874998765, 0.0143199537928174, 0.301901965406671, 
    0.0353913631743256, -0.05044211867069, -0.0429000143604159, 
    0.207957021076746, 0.278391703706137, 0.363403136267624, 
    0.110458252991245, -0.47993095073395, 0.532376538703858, 
    0.529903233564374, 0.193330506311756, 0.261936861580194, 
    -0.309912352804319, 0.802401428777971, 0.281032965338549, 
    -0.127902332273793, 0.327811783594404, 0.21807606988458, 
    -0.110762280198413, -0.190136368201005, -0.0151110314555579, 
    0.447855101848784, 0.142391143035057, -0.394166325017213, 
    0.0398554470176241, -0.358584279615821, 0.0411337376008829, 
    -0.322001102576507, -0.0114292397361539, -0.32539413723673, 
    -0.0282712500211397, -0.452191710754769, -0.179600796297584, 
    -0.141038143533035, -0.319189243973978, -0.033790958140981, 
    0.012818421230707, -0.0179067100271319, 0.000817009071458999, 
    -0.0089644534235927, 0.0109422694769398, -0.00976837732674837, 
    0.0218931033162901, -0.030712979837106, 0.0827236972896881, 
    0.33881119508304, -0.119510709599661, 0.333985507910627, 
    0.431803190995805, 0.0682009213515488, -0.0656371279099744, 
    0.305536263447685, 0.573230466309545, 0.481498040536049, 
    0.238859420438541, -0.0203656229466725, 0.610674925336629, 
    0.247418639847303, 0.0138589355613084, 0.0378266351529968, 
    0.442454308033574, 0.120599216376708, 0.164704644080199, 
    0.674372655269914, 0.1928462005076, -0.0172057845999879, 
    -0.00362149961154362, 0.0209904782896609, 0.0054567213524412, 
    0.0167677404120939, -0.00163837708296422, -0.00135535969484092, 
    0.0285619406447341, 0.020580890203841, 0.00682169971585052, 
    0.17641746727253, 0.0606126163457563, -0.133786977017956, 
    0.115903647745509, 0.488385502277849, 0.142053762674754, 
    0.00959616490905139, 0.0747854193724861, -0.113256324715875, 
    0.601510461197351, 0.201219691192291, -0.04484370934647, 
    -0.0893305936119089, -0.109623530346512, 0.768386723376254, 
    0.299050295848868, 0.102416661406432, -0.177760133233639, 
    0.589900561622818, 0.120006183843974, -0.0719389548241037, 
    0.0999932577246491, -0.181525240033367, 0.0499912139693969, 
    -0.277722868465088, -0.0859198765298826, -0.0952396359615737, 
    -0.172053239741793, 0.0446628711131637, -0.18337258243229, 
    -0.00227604646016862, 0.110803553334849, 0.146602733881122, 
    0.16094705861029, 0.226373115201613, 0.243546291700099, 
    0.188329295990344, 0.138127891602626, 0.186633707668324, 
    0.27706906449327, 0.25804598710721, 0.198953161003726, 0.164226501906446, 
    0.166803783712764, 0.177813909274928, 0.156060713243797, 
    0.156941798429402, 0.209002490036245, 0.185387612259109, 
    0.131034274335094, 0.195992111076872, 0.187726675813578, 
    0.111336923747245, 0.305581440814271, 0.284979999175551, 
    0.0423193781276771, 0.228434443896798, 0.452211479453016, 
    0.0906077661325455, -0.0179509431777854, 0.108907660002449, 
    0.565020211637504, -0.0630375924167307, -0.248726803797619, 
    0.171080453576277, 0.354375281150723, -0.0727717790553044, 
    -0.337577449480042, 0.320825570330976, 0.0759536943541698, 
    -0.322219645089892, -0.165264579743271, -0.0013004767090322, 
    -0.245931437980627, -0.116001281662379, -0.130997908998809, 
    -0.0501486184243923, -0.3079530030171, -0.200776662102292, 
    -0.248710738129077, -0.235511491355318, -0.242491545013145, 
    -0.114314860095888, -0.236553261346706, -0.0519728382788465, 
    -0.200507861718755, 0.0121607282190516, -0.000555120321118319, 
    0.167028005886291, -0.358533286419423, 0.0433634606780425, 
    0.0446514391362551, -0.0276698471198235, 0.0693295096245493, 
    0.236024158721105, 0.184128512452727, 0.103317459559315, 
    0.0835030790309554, 0.0903404236515419, 0.0696641501835734, 
    0.178235330193768, 0.301939072928765, 0.392531857842211, 
    0.29763979262593, 0.141163528919715, 0.265370635677955, 
    0.517113407924971, 0.269813079327215, 0.0813884977145695, 
    0.260350371822498, 0.186625379581291, 0.0601144793511667, 
    0.774778431639888, 0.414407998492747, 0.0661685704872631, 
    0.142681780398344, 0.679165753285392, 0.0241177824151494, 
    -0.0980680194999862, 0.178565114091684,
  -0.145824049230911, 0.258883920113271, -0.413717577000656, 
    -0.0163722117377654, -0.468627778231157, -0.3779033361142, 
    0.133793526097864, -0.0931284870573453, 0.24940711308041, 
    -0.449383640681589, 0.0290980381402999, 0.0322705496241927, 
    -0.0331803782205542, 0.0620636247173782, 0.0105632307812296, 
    0.00386691462384482, 0.102256120669447, 0.0679615484865612, 
    0.0400589399188346, -0.0914932919631237, 0.0307802773735599, 
    -0.0683370272438474, -0.025703616811575, -0.0618890597143517, 
    -0.0285412443271633, -0.0397363127752681, -0.0411058837929709, 
    -0.0224019908690413, 0.0399540228023016, -0.113668760773838, 
    0.0686307664053529, -0.0263666984241178, 0.301316806287459, 
    0.222418435612088, 0.162133588383162, 0.237946651487014, 
    -0.089257476354493, 0.486585809720983, 0.232849345280158, 
    0.131843322334021, -0.387678073853464, 0.241723691540471, 
    0.398912797388191, 0.13189745438465, 1.02833504950405, 0.592813270272116, 
    0.0723033502143559, 0.181866523311109, 1.03370856603282, 
    -0.0750701289296466, -0.12653046798327, -0.0282111615373359, 
    -0.0202721535282454, -0.0505046743696795, -0.20453171228435, 
    0.0882852314560995, -0.0333838110298157, -0.0711505684519603, 
    -0.105905295923264, -0.0506243428797357, -0.10383712635401, 
    -0.0993482586337293, -0.106172620846477, -0.0258543856639621, 
    -0.12562962509079, -0.0203956352915281, -0.149634751662529, 
    -0.0523879953603348, -0.0793401174384279, -0.0635737782526515, 
    -0.00719280533429469, 0.0637572436426252, -0.00731685620970148, 
    0.00777749134967602, 0.0489559452756322, 0.0172351308065547, 
    0.0316868988529027, 0.0720789864667306, 0.0865369849185514, 
    -0.0576823442912025, 0.108831546062679, 0.2383597302574, 
    0.107137242846085, -0.0141938075024029, 0.232146386903538, 
    0.3857561651835, 0.254839317093866, -0.0663977338236289, 
    0.56876501967479, 0.141705594395738, -0.221466303977542, 0.3861301440649, 
    0.413153435572016, -0.00742294868438689, 0.0562038662182728, 
    -0.11004887580222, -0.031275277989689, 0.268372295608762, 
    0.0054471466113275, 0.819551829930598, 0.841387719541873, 
    0.0391525209543554, -0.132443245853055, -0.120711973623656, 
    0.157713897482137, -0.170124743035426, 0.202900554074428, 
    0.199172407162036, -0.106192180801148, -0.0759958879251891, 
    -0.000541105016978252, -0.180510301025621, 0.0940809883748878, 
    -0.066553249308543, 0.119437102956308, -0.152480169583186, 
    0.158291872161542, -0.275074200069613, 0.101286555094172, 
    -0.152255703963857, 0.235760758654843, 0.033715415769544, 
    0.0538775500557945, 0.137355988720251, 0.199475277757202, 
    0.450566495763062, 0.335634337153066, 0.033322576165131, 
    0.00150378035606558, -0.397369680081138, 0.0677091863229278, 
    0.657183375407411, 0.136490560118121, -0.181275795620816, 
    0.0780671379910826, 0.531865916456464, 0.205522433649341, 
    -0.0938581139270013, 0.382398152493885, 0.389511633277625, 
    0.0577402658507686, 0.0321705685993073, -0.00559464850251572, 
    0.0193678594852117, -0.00774905893736243, 0.00739163154687672, 
    -0.0196215618432314, -0.00587236619205711, 0.00999488845479715, 
    0.00819821044206448, 0.0518824304031072, 0.0862946346054284, 
    0.023717878290549, 0.292877453627439, 0.350835555952568, 
    0.134151573704681, -0.0531793124118985, 0.559341957001545, 
    0.120403566128939, -0.306690617591847, 0.10044640606387, 
    0.628210860490434, 0.262238114883385, 0.166678818705565, 
    -0.0560629972578285, 0.344201796085743, 0.304284442719395, 
    0.410028531408841, 1.34495896650458, 0.101346129576804, 
    -0.362398881514617, -0.173305439747531, -0.0494206354452565, 
    -0.200025362197113, -0.0135284127110958, -0.190845670867215, 
    -0.0854855392452451, -0.0613298517557683, -0.196227671116902, 
    -0.146437428650407, -0.0116101725899069, -0.0184012726778412, 
    0.0863472959565253, 0.0575460836484179, 0.123922519217586, 
    -0.179714735962005, 0.100234337993349, -0.137326245555321, 
    0.0149000518167137, -0.112956232369905, -0.00961583752958993, 
    0.028398105861276, 0.0371241974126962, 0.0395888550234205, 
    0.044343195713158, 0.0628591873354029, -0.0610766691075972, 
    0.210585517975626, 0.0657022629066672, -0.189940658948496, 
    -0.0849752224673942, 0.425773356381562, 0.180945045079386, 
    -0.118429007453956, 0.444089778180371, 0.497906329858521, 
    0.14161716668527, -0.162895017818884, 0.132009857825155, 
    0.276504927649799, 0.206129121597795, 0.696305674234443, 
    0.311218891775375, -0.0456010970542326, 0.087065309013028, 
    0.141862187710017, 0.0613200540422168, 0.947642600806164, 
    0.284432975544564, -0.0475012670599785, -0.202449747087369, 
    -0.0101641461217399, -0.396762452535737, -0.185571495580903, 
    0.0630862707969023, -0.262251209447653, 0.0628496659760341, 
    -0.0880227031050265, 0.0146022669225796, -0.30532430619344, 
    -0.0479134704805725, 0.121098900982794, 0.158887411748984, 
    0.124078002763485, 0.226131514548043, 0.372010611642876, 
    0.300639371877242, 0.168697169933135, 0.145993776561908, 
    0.297034518671854, 0.371050832813841, 0.31158635322789, 
    0.258393743449319, 0.261367383026253, 0.261841476123947, 
    0.199011060291071, 0.203452945290023, 0.349668825910708, 
    0.224187153839713, -0.0346887361759573, 0.206166382186999, 
    0.468707969953435, 0.227742499258721, 0.104135402316564, 
    0.190558464271237, 0.0912696613326618, -0.0259452513307558, 
    0.623222779259356, 0.493354545157373, 0.0457127465948819, 
    -0.1794946609888, 0.0477263556657303, -0.327533143564844, 
    0.69741524579122, 0.921682148615236, 0.302287928070736, 
    -0.510935954990984, 0.593114063800976, 0.445865497898162, 
    0.0209960830395427, -0.24451286204297, -0.0540299417512185, 
    -0.168481373040682, -0.133753911040599, -0.104799696032549, 
    -0.151007595640386, -0.0663966171636053, -0.135984186347977, 
    -0.0218926222870328, -0.157496228279011, 0.0384398042742123, 
    0.115958009929307, 0.157831014513412, 0.17692034522211, 
    0.172474503967547, 0.163974799064223, 0.156383405009169, 
    0.171817860520911, 0.186577273929124, 0.177474206419995, 
    0.184610066878717, 0.182474282082407, 0.184400503557792, 
    0.223013235839154, 0.228007093898039, 0.152950061675556, 
    0.162925437718954, 0.342958486768993, 0.19992283124379, 
    -0.0199216279044553, 0.068386021581416, 0.505530822857433, 
    0.188428246768551, -0.0532844291688181, 0.0712052992176225, 
    0.369565742514674, 0.276162625308821, 0.429667822719214, 
    0.372750636210399, -0.00943025617966427, -0.139257537107003, 
    0.874563642277675, 0.421907675352881, 0.0655308643282515, 
    -0.0911583736302705, -0.320856301887398, 0.443011001027399, 
    0.395929320697417, 0.184722002638383, 0.521183794761532, 
    0.478020709820022, 0.320614106532043, 0.126851184361478, 
    -0.1470730055595, 0.203057490616524, 0.218419931592411, 
    -0.119940725941142, 0.138958866730933, 0.410973931423783, 
    -0.112764162599229, -0.0555961616114696, -0.0180483689061136, 
    -0.0438883060156877, -0.0252026562683772, -0.0424282533936526, 
    -0.0184646786150325, -0.0418710398141781, -0.0153079816992328, 
    -0.000935280199467814, 0.0233479606697633, 0.155046891068672, 
    -0.113637588981869, 0.255005358858364, 0.273738567499481, 
    0.146667285936333, 0.352969628723371, 0.276565110680933, 
    0.0351442499782662, 0.691044172962139, 0.240135515545414, 
    -0.155129781409851, 0.182550264289864, 0.548898880456609, 
    0.310570465707065, 0.121533812097641, -0.327373497291624, 
    -0.118499614108074, 0.596914130818276, 0.228492070280839, 
    0.243313613286277,
  0.0840294844403773, 0.169026562407678, 0.160688274533854, 
    0.317058323007232, 0.214815150153585, -0.0771452695509581, 
    0.177396837806354, 0.416541758463446, 0.36833890531061, 
    0.406761888671143, -0.135401647985955, 0.509638879161287, 
    0.439316532311655, -0.0860679400418376, 0.414892560070924, 
    0.705254863035063, 0.199807616231142, 0.320904241748235, 
    0.0772073728970368, -0.618146642430024, -0.469873072355995, 
    -0.00730115751701604, -0.203829338129188, -0.182144577365221, 
    -0.148184460980809, -0.148106743285917, -0.0407612615603842, 
    -0.203513440338643, 0.168055673084756, -0.247386835694064, 
    0.151161919766289, -0.00963429415642994, 0.116088907888804, 
    0.0450097958056146, 0.174017413104172, -0.014984243826763, 
    0.137387387107793, -0.0209587621193378, 0.101926844822788, 
    -0.0617974007978481, 0.0237122726882853, -0.0793726301957619, 
    -0.0213775577661475, -0.0830704880690598, -0.0460806435859429, 
    -0.0586432824527127, -0.0529681009594795, -0.0341755768796831, 
    0.0944058681406459, -0.133211172316657, 0.427514864899167, 
    0.158998439035692, -0.236356490108655, 0.178934676025088, 
    0.42815834264409, 0.166623256829523, 0.0478364293186681, 
    0.533432693151693, 0.3389586194553, 0.0978143667907562, 
    -0.101505415594046, 0.156929992250954, 0.239823146873274, 
    0.29688978281459, 0.298238655407572, 0.111655147579703, 
    -0.0108114098207523, 0.293152740956384, 0.117019082519843, 
    -0.0138908322308255, -0.0462171222293221, -0.22830203685579, 
    0.106082863721394, -0.122839711705295, 0.0756660873963813, 
    -0.212552618853168, 0.0554098047940841, -0.125315457479394, 
    0.0684067966364974, -0.348545251744307, -0.00573215060467767, 
    -0.0855527893917235, -0.0732446074930804, -0.0735923428789246, 
    -0.0635410101045036, -0.0696569241922664, -0.0570356429202942, 
    -0.0340730732617853, 0.208308540105296, -0.178761949963835, 
    0.393632125408869, 0.286492559813352, 0.557216371287438, 
    0.351927547167916, -0.280305760401971, -0.0209408095060996, 
    0.600410978891454, 0.365289505821187, 0.171698372852761, 
    0.0138341063367755, -0.0349621280429066, 0.311785466891171, 
    0.254782399037731, 0.142142980001567, 0.109083904490559, 
    0.101804510711849, 0.0985665825047049, 0.114287525845367, 
    0.137068148221078, 0.112892360164204, 0.0320265013218372, 
    0.0300885969718862, -0.0246833626690015, 0.0151034230570211, 
    0.000691674587748187, -0.0203288096320528, 0.00347031111773784, 
    0.0415774259784961, 0.0381277663740864, -0.0156171227059118, 
    0.0195483676263515, 0.0347810393044417, 0.122037679988138, 
    0.352496109603176, 0.205341466927681, 0.060692910892815, 
    0.298157204467073, -0.0777674930907604, -0.314277708952663, 
    0.00351987525721298, -0.368684883967975, 0.380238583621068, 
    0.507586981554884, 0.141627611265159, -0.0739525459144494, 
    -0.486789781465112, 0.510434720341527, 0.525867563679644, 
    0.246385203603064, 0.0815432822910696, 0.0672540220720359, 
    0.276767709089993, 0.0979303096012988, 0.0109175859629269, 
    -0.00908666048617233, -0.039022176754991, 0.0231381137716413, 
    0.0574846655903777, 0.0181973205657038, -0.0132359534875026, 
    0.0251402252509813, 0.109044381811205, 0.0953087795199232, 
    0.0580445732696919, 0.0660738210907231, 0.101514339275982, 
    0.0715622005052, 0.0532189495021977, 0.100611477272042, 
    0.0747135046405974, 0.0445077854787145, -0.0122717627972033, 
    0.366396141376989, 0.264506614543185, 0.0825268312705739, 
    -0.0855364655489719, 0.0429561222025941, 0.349589945589707, 
    0.257851359161391, 0.159132207291513, 0.271403072423572, 
    0.276487224325555, 0.115595171086912, -0.00899690256755305, 
    0.242544072775083, 0.540347174022785, 0.476712178865388, 
    0.182217282206718, -0.143386111750432, 0.129920508299697, 
    0.679096750351482, 0.072175334499526, -0.0592126879977526, 
    -0.177820040829268, 0.214540030093558, 0.593326501385013, 
    0.238685592428856, -0.084285933064043, 0.300005157003005, 
    0.37551253612169, 0.0600289583077763, -0.0571017528375335, 
    0.136151885920597, 0.274923777517533, 0.0381589618691221, 
    0.00932421476525799, -0.297851135783752, 0.00583311753708797, 
    0.392077052537682, 0.0836784499331514, -0.0440184639161235, 
    0.0411543131325265, -0.179927521822288, -0.00103989478660534, 
    -0.119770204896368, 0.0322134419922738, -0.197807564699585, 
    0.088417941788262, -0.174911480964709, 0.0504857022904782, 
    -0.0910317464513642, 0.0386335702949375, 0.307627827444152, 
    0.108058957540683, -0.0420752158688523, -0.0674504546752904, 
    0.169245897545026, 0.569989160824231, -0.146107799378707, 
    -0.17591035725275, -0.320029032711242, 0.411068781423603, 
    0.517164166755206, 0.142519983660275, -0.321869689503054, 
    -0.0666258675842921, 0.690895746120384, 0.153344536296973, 
    0.54509663512622, 0.999434987776382, 0.0116904783700621, 
    -0.0371319057065854, -0.0321633023604914, -0.0649368000433434, 
    0.0988800860409216, -0.111218098154109, 0.216203945827307, 
    0.379025362910134, -0.160140111650542, -0.150778396908459, 
    -0.089758683940257, -0.169851621835546, -0.0445136927045079, 
    -0.167183598572442, -0.0948309029745359, -0.254977789801952, 
    -0.140133269819862, -0.138717338193415, -0.140474364307678, 
    -0.165436533524038, 0.0419678589118669, -0.0654286713440477, 
    0.0807332469318387, -0.0505106824899669, 0.0255743130288539, 
    -0.103507192121643, -0.00352704558130071, -0.0329975023017271, 
    0.042410299186475, -0.173357500302608, 0.00754480873546969, 
    0.0485496177995308, 0.0703381820704876, 0.129534149915291, 
    0.112812410248192, 0.0306449836063981, 0.0471358564064661, 
    0.349272990502657, 0.229474531102496, -0.224056108758315, 
    0.509518586034784, 0.316960655773992, -0.104758968359657, 
    0.194465306874081, 0.68415270823825, -0.0401767886470629, 
    -0.0238997243913288, -0.0629912965952944, -0.207787114383811, 
    0.901278698069621, 0.108655982852732, 0.0646208944170776, 
    -0.37551734333261, 0.677066932248242, 0.414201383920171, 
    -0.373966034078343, 0.55854500118159, 0.504820832850017, 
    -0.1262796249941, -0.0590241115052121, -0.298042357999733, 
    -0.282685487299833, -0.179957117478731, -0.280452402022371, 
    -0.179256503956857, -0.263372177062266, -0.0915499878740896, 
    -0.260904519742094, 0.0239833248247306, -0.28545051421663, 
    -0.00453459950526862, 0.098480634425856, 0.124562167944152, 
    0.134787488736913, 0.138134292579225, 0.116557772129598, 
    0.107920412852379, 0.202090296182149, 0.160376729908487, 
    -0.0397306995860296, 0.212318641424426, 0.370905397445457, 
    0.137349622357294, -0.0259605268550879, 0.434579322881601, 
    0.381154935826187, 0.227569778632483, 0.208229553943757, 
    0.198124604584714, -0.25961815211651, 0.551657374087341, 
    0.452343959707876, 0.143395893092038, 0.0870675861751509, 
    0.00781977766528393, 0.729878961118687, 0.0671823316638866, 
    0.0630131672595692, -0.0623633840909121, 0.605966264007005, 
    0.0620787809660704, -0.169101032590241, 0.34433210524631, 
    0.328176492036646, 0.063665542275472, -0.00994255704246379, 
    0.024519402436283, -0.229653446435548, 0.146078870700806, 
    0.140384211757499, -0.227989325261393, -0.115307120079419, 
    -0.199112262475843, -0.0761787553027984, -0.175973469567382, 
    -0.131255608076896, 0.0561180001886233, -0.19328145232224, 
    0.0941634759017603, -0.140449669434536, 0.0870262231046914, 
    -0.0315922042070145, 0.0417394131670717, -0.00453665468254337, 
    0.0399286560476229, -0.0311852476703079, 0.00388511510058362, 
    0.0625332648491679, 0.106814868527658, -0.0765369780357987,
  0.57954382553973, 0.222888592142458, -0.0258994478725558, 
    -0.112507864731029, -0.182942386063532, -0.0261529584890477, 
    -0.137963331648937, -0.205382725165485, 0.0561941881208946, 
    0.012222512434838, -0.0315872307948843, 0.0647399052765783, 
    -0.100289447797207, 0.0350304936452232, -0.0136228806298219, 
    0.0499923639232712, -0.192793995950438, 0.000229623472167234, 
    -0.265715072340249, -0.154970774576104, -0.0166435693699044, 
    0.064020849002043, 0.0898809728660669, 0.0679938423430322, 
    0.0706034155305411, 0.0963541990341955, 0.113900584575936, 
    0.110677014065511, 0.0931462590924717, 0.0540100376390664, 
    0.136877484309043, 0.154262213643479, 0.128828133965822, 
    0.214223045758472, 0.307867531158863, 0.194909432062279, 
    0.0662201331253813, 0.183703968635962, 0.349587225773515, 
    0.353468243195034, 0.184412826132846, -0.169235065070555, 
    0.095357718344533, 0.472098123656062, 0.2538760580689, 0.160156339153292, 
    -0.19747088179959, 0.249576430238643, 0.397051148334051, 
    0.206572893518986, 0.0222271608432333, -0.091825325640137, 
    -0.0656876839074701, 0.46246033527034, 0.0357335358444254, 
    -0.0157412304621168, 0.0407219651546676, 0.501588658911222, 
    -0.0341757085485582, -0.0491458277760888, -0.141143126114793, 
    -0.219831557363903, 0.129495236964717, -0.341179663023603, 
    0.00225677309511971, -0.299428642909298, -0.160966007047294, 
    -0.149375065946626, -0.151216185656294, -0.147293994992454, 
    -0.0220764715567603, 0.0857201426002271, 0.105500889958472, 
    0.121921537850132, 0.158204966925472, 0.143175407836708, 
    0.111986399846528, 0.136097413147464, 0.0972093974000037, 
    0.0314235764939855, 0.182200259001872, 0.21730764367249, 
    0.0971713816139082, 0.0514159741593353, 0.304677557423693, 
    0.379926830266527, 0.197303242973165, 0.0646212800814751, 
    0.035432431350393, -0.114549750698218, 0.637475120324665, 
    0.294693496943693, -0.0459246716665252, 0.278745665042589, 
    0.389753846751856, 0.0679052358191018, 0.391419851829509, 
    0.546597121737731, 0.25805167529045, 0.34950403275245, 0.350602939138217, 
    0.051001469672916, -0.0300599081222273, -0.0242160868900831, 
    -0.0831280018691238, -0.0015426389484922, -0.132319603093386, 
    -0.181885502647905, -0.00175926245484243, -0.0551712982786805, 
    0.0894608478086242, -0.140626046935749, 0.0783942765372995, 
    -0.0813357886235943, 0.0544496193484519, -0.186190174595896, 
    0.058241066126583, -0.124170689743493, 0.0422055392974051, 
    -0.268776012503077, -0.0374845211414563, 0.0239490562032894, 
    0.0392196630056957, 0.0835152158035152, 0.100813926159058, 
    0.0581246754553182, 0.0633222559876345, 0.177684201507967, 
    0.0787609995813573, -0.129849468551775, 0.0526274647920299, 
    0.396116658911663, 0.192834933909517, 0.0411918889323525, 
    -0.12042902262591, 0.32611517443794, 0.690596960490375, 
    0.0644931008925948, -0.268062074313143, 0.0548055103008446, 
    0.597289178855091, 0.0632130377526403, 0.192899205758867, 
    -0.401066732649889, 0.514253360221499, 0.496195970629419, 
    0.143141894931755, -0.214428963750982, 0.0817438922647554, 
    0.472153818370163, 0.21777760723376, 0.192042792991946, 
    0.114480042760426, 0.0588451772577095, 0.0505963803878665, 
    -0.06605215258443, 0.113607873354323, -0.222184265262011, 
    -0.21473399054593, -0.159603480193561, -0.093054791270112, 
    -0.287519560131873, -0.107505627438033, -0.0805170091850417, 
    -0.206748376869143, 0.104236523147628, -0.1860353997239, 
    0.0500775068389137, -0.216656162699583, -0.0585706056985118, 
    -0.0293416846944389, 0.0357873927193115, -0.0067055064522713, 
    -0.00533704172505078, -0.0268336504392853, -0.0253133648672168, 
    0.0483256969646454, 0.0185135415017562, 0.0903436298250828, 
    0.0211859434966486, 0.0806633294294936, 0.0829070467046415, 
    0.0777525335440054, 0.0912197261930921, 0.095510535228377, 
    0.0735208451211607, 0.0681568225260615, 0.122313044900288, 
    0.0976407080412683, 0.0249031059525337, -0.0246813369864128, 
    0.243034852556147, 0.265498379833439, 0.087546663281461, 
    0.038198842495444, 0.42255146337893, 0.219435210352268, 
    -0.0300193586262762, 0.0851697733947174, 0.54456274178837, 
    0.169534182628016, -0.0930143974487812, -0.0234435980363297, 
    0.475161435693731, 0.192076070980074, 0.685633993106668, 
    0.503414897895007, -0.261882916705592, 0.31012542056318, 
    0.512785804704561, -0.177741892701271, -0.0877973859851608, 
    -0.0204226211599905, 0.0075977257373625, -0.183669290396281, 
    -0.190685811607468, -0.00377905273008662, -0.128868592539764, 
    -0.222273275107802, -0.104932582752262, -0.149119412869455, 
    -0.244600151072524, 0.0265061582589925, -0.00662599646235006, 
    0.0976063936251411, -0.175418568135983, 0.0602128447554069, 
    -0.128420551942976, 0.0373488078002827, -0.257505287093002, 
    -0.047304533984052, 0.0400970370522935, 0.0380003028576884, 
    0.0397226462084756, 0.0920238955697232, 0.142043157082731, 
    0.134540207186291, 0.0855546016915932, 0.0991750745656496, 
    -0.200395318007862, 0.460256106041364, 0.278327761407239, 
    0.0804596521781329, -0.082744092913432, -0.00135598087980487, 
    0.0315080751999629, 0.75465301907739, 0.446440275026181, 
    0.241533503989825, 0.620588793545915, 0.121936871757026, 
    -0.141850179792946, 0.214316332268323, 0.374839378332827, 
    -0.191562817525437, 0.177591450686153, -0.00540962980269725, 
    0.999120710668004, -0.0170739814897369, -0.32323258331927, 
    -0.318490473417821, -0.0725438282729063, -0.209304141934544, 
    -0.165462520868343, -0.166203006295638, -0.171509265100286, 
    -0.0999680371786396, -0.182954363758262, -0.00580212968434379, 
    -0.210512052165405, 0.00713120444064919, 0.100710306947809, 
    0.132303470103564, 0.182685815350707, 0.257207087825257, 
    0.235750252125032, 0.164087460497565, 0.139390047413229, 
    0.232745674133159, 0.365925362320648, 0.300483556857484, 
    0.110546767031284, -0.156537545010826, 0.272607606784426, 
    0.540809461687963, 0.184060248172173, -0.0431498440691429, 
    0.169024574026469, 0.392071452247183, 0.0545825579415529, 
    0.348006721974246, 0.657542761210343, 0.0611527020042489, 
    -0.000887372943050205, -0.200855398971969, 0.47238777613492, 
    0.321907720961325, 0.0692076800140877, -0.0561529769759215, 
    -0.107077023577455, 0.526139774118962, 0.128189868780041, 
    0.0179552605556038, -0.0442274920715642, 0.100020167543083, 
    0.213847183551263, 0.378966710892037, 0.338917220070274, 
    0.202194697276575, 0.198977417402878, 0.251725715489539, 
    0.368679539858113, 0.242709961454261, 0.0495206146546333, 
    0.341039145548075, 0.400795717504485, 0.0976131469042498, 
    0.0236814541746096, -0.0754492474136681, -0.192612501094825, 
    -0.210464983019153, -0.206184076263369, 0.122452377099573, 
    -0.148087686486876, 0.0947954206502485, -0.0515325078555674, 
    0.0611255550722377, -0.101517256848751, 0.0399105013411057, 
    -0.237672696127319, -0.0240211410743947, 0.0323250659346321, 
    0.10891061533711, 0.168450063598336, 0.138412045810543, 
    0.0852926532636313, 0.0690478147373744, 0.170073650653605, 
    0.163354872161083, 0.0593966490987964, 0.0567698423070673, 
    0.256819234788784, 0.298170535748104, 0.187535504990961, 
    0.296037062484737, 0.401974392024691, 0.198046615646233, 
    -0.0226088778268554, 0.277174842611428, 0.676473648687832, 
    0.256326544064321, -0.247250521289355, 0.409734202861841, 
    0.555886980460549, -0.110325204785824, -0.117354719346964, 
    -0.0114068667348409, 0.0686970560172093, -0.0818927773838824, 
    0.51452445230069,
  -0.0504914896159339, -0.251234894863309, 0.0798772585604767, 
    -0.176564602008132, -0.00829949212030555, -0.175908514965137, 
    0.00273992875477688, -0.129867694474259, 0.0695975853220683, 
    -0.245178647046093, 0.118194746820297, -0.0431976791320749, 
    0.179273337866212, 0.394135072955231, 0.144995496029391, 
    0.030493279784658, -0.216291074362745, 0.346029147938418, 
    0.461589647398339, 0.120491253392298, -0.0439172642813584, 
    -0.0447132646202192, 0.686996968682671, 0.27629835948693, 
    -0.247468943963639, 0.351875475528624, 0.794315822045696, 
    0.213048223873874, -0.169111530744187, 0.497296115717616, 
    0.491372315623926, 0.133692889790468, 0.0329669889802541, 
    -0.168059723740861, 0.169935511673877, 0.626036518325721, 
    0.122818415338078, -0.180236352997199, 0.139534734925923, 
    0.426710668563556, 0.066075637006563, -0.0580856611070449, 
    0.178265990231731, 0.336891617598931, -0.132816160285995, 
    0.158183262886197, 0.471952765512676, 0.169470173604651, 
    0.0485775787786646, -0.0322836764709986, 0.0806067353957461, 
    -0.236389638639736, 0.215543061406845, -0.12642527913652, 
    0.053554308089491, -0.173090627298085, 0.00661175627986078, 
    -0.138843421208448, 0.00205098166811518, -0.291611543751256, 
    -0.0305553054238975, 0.0377150307784914, 0.14592192348825, 
    0.173153544829587, 0.140663716650617, 0.0774234755048744, 
    0.0729988334393591, 0.159929790913081, 0.13611601063859, 
    0.0670658771889877, 0.0489205623660144, -0.0250262489955206, 
    0.0135609872375341, 0.00647227449864701, 0.00672737364682395, 
    0.0136138605333428, 0.00363305076833789, 0.0363391103655055, 
    0.0533107669730147, -0.0675258540397524, -0.113911626653899, 
    0.243560490628025, 0.357490333107907, 0.364440506332293, 
    0.236063274490826, -0.0286521036740914, -0.256129356419218, 
    -0.195610402555556, 0.723150045186344, 0.0997937564963776, 
    -0.104049337575925, 0.127548675151682, 0.253860466514148, 
    0.0554415575985479, 0.45532784097255, 0.354367697722097, 
    0.0552367312437274, 0.392414002075474, 0.414428137703904, 
    -0.00187264001761481, -0.0789734978997803, -0.0889472921821531, 
    0.0111602784329725, -0.0815823563885881, 0.0144680886902193, 
    -0.101073385301605, 0.00596798909230185, -0.0414364715238423, 
    0.075369732303823, -0.0600513995811136, 0.204531730752768, 
    0.0187514130313371, 0.00539860364441917, 0.417440498418294, 
    0.235697239584552, 0.137929326620278, -0.0931821451454264, 
    0.340784774853782, 0.220895636408272, 0.0174133411795766, 
    0.0020215210217955, 0.70449153073912, 0.431377615095409, 
    -0.231646909071825, 0.791833235721024, 0.385849288272903, 
    -0.120061378158536, 0.592973704551457, 0.576492219689001, 
    0.04790112760673, -0.0875507304516037, -0.0885184079609066, 
    0.0388525989260662, 0.0166977163808128, 0.0646142714443582, 
    -0.0782704233839936, 0.0185061140799457, -0.000584320461444618, 
    0.0386493262172444, -0.093064038591385, 0.0190447901576811, 
    0.0663735004115202, 0.163149477543605, 0.304869958530808, 
    0.358022208987645, 0.164434094921851, -0.0445205434912268, 
    -0.123683763683863, 0.439097779484906, 0.565830838435845, 
    0.295864623250431, -0.169463096691249, 0.560667249795406, 
    0.486895985122086, 0.15208082691334, -0.0659539955113607, 
    0.72565993724818, 0.431820155907047, 0.217631587108318, 
    -0.187038167816333, 0.418405142405793, 0.410748966314422, 
    0.135341374643532, 0.11256664273109, -0.270722048283827, 
    0.490785176705656, 0.286144032476676, -0.0792386569619266, 
    0.285987305492734, 0.610047760115363, -0.107870899702698, 
    -0.0415047339750275, -0.0714600305681085, 0.0193036873368218, 
    -0.182478153754654, 0.0996040731890587, -0.180752797502368, 
    0.427003173836003, 0.446585848757072, -0.193433280099321, 
    -0.248471583716244, -0.0841598587347885, -0.175341144142249, 
    -0.137594622831629, -0.170333185085181, -0.153381344827125, 
    -0.113061266344775, -0.1627691198441, -0.0373939292712855, 
    -0.172167321694184, -0.00996335555372824, 0.0655180981033658, 
    0.0770210298032935, 0.0871086226429564, 0.102318267323241, 
    0.0903540720581093, 0.0315780961755109, 0.0293841189095484, 
    0.203998019291648, 0.181550942373178, -0.0674004830862188, 
    0.356558830621928, 0.412803246891482, 0.175242260179387, 
    0.281767038238057, 0.401533600731884, -0.0362336251890497, 
    0.540608938386475, 0.598287635524815, 0.0717206526195787, 
    0.402187558016887, 0.729259900532158, -0.0250580128914111, 
    -0.186174848125382, 0.0236427585904659, 0.515508408454996, 
    0.190303711896265, 0.331457358593426, 0.245120556558717, 
    -0.226920067767291, -0.293028091695931, 0.146364091758734, 
    -0.376187774246545, -0.161521099206756, -0.0346406436179961, 
    -0.204324618088307, 0.0285824127627359, -0.113408742772182, 
    0.0489650044489451, -0.227427805436807, -0.0406102433635196, 
    0.144321692806875, 0.213297190159053, 0.0960403467291379, 
    0.185896303973006, 0.498473577064165, 0.29444628368865, 
    0.0463176579440695, 0.165350744604338, 0.483593328154547, 
    0.343654343699817, 0.21783900718203, 0.181804268266113, 0.15505638835718, 
    0.139952362690895, 0.175279303059384, 0.191017055001652, 
    0.192130076226973, 0.209024461302055, 0.177978717132288, 
    0.129518938663668, 0.114290949873315, 0.132043637026479, 
    0.206308258269757, 0.192068706170233, 0.0859035364338766, 
    0.120863375490645, 0.379816186123675, 0.17483581982515, 
    -0.11875413333634, 0.286423805745307, 0.36453994775441, 
    0.0190328025388921, 0.102090437907033, 0.644136520438216, 
    0.160692209342443, -0.197279002046204, 0.270908222003743, 
    0.498283684314876, 0.0308943443050494, -0.0114717263509509, 
    -0.270652077321789, 0.354915218903507, 0.366019086336968, 
    0.127720999947967, 0.0875600522563425, -0.05122531173034, 
    0.628802173636616, 0.114780187508028, -0.0146842149936571, 
    -0.386614086133285, -0.0492302324006392, -0.257800618050758, 
    -0.241917302292716, 0.0691788877105892, -0.250946809734147, 
    0.109141645584036, -0.154411587349019, 0.121610913546978, 
    -0.252196617992198, 0.0312895662295202, 0.0811446046206821, 
    0.128670361048644, 0.121291502298577, 0.125399435959642, 
    0.0689959191554707, 0.100541508046337, 0.126726024868837, 
    0.0874401414861078, 0.0047029571340472, 0.0335363124105339, 
    0.0069499650367877, 0.0152875433894985, 0.011159094412637, 
    0.0198800822182583, 0.0201856602232737, 0.0370656613687507, 
    0.0678807233166017, -0.201746116021352, 0.127156609046593, 
    0.373361623941716, 0.0491997571115923, -0.357599737172968, 
    0.239606512924799, 0.333930005782862, 0.611859365549302, 
    0.450155326516153, -0.113582438920508, 0.508701432038466, 
    0.519270069730755, 0.0696871766426137, -0.0184016063568349, 
    -0.14004197936082, 0.152684644021835, 0.130868396600987, 
    1.02471786311758, 0.5475177428984, -0.0114714118232651, 
    0.574158945936687, 0.441490961590744, -0.193634510814693, 
    -0.0452843186392846, -0.0707832138285169, -0.0399963193605821, 
    -0.068056237173917, -0.0004915205773766, -0.091700528835146, 
    -0.0121450953080058, -0.058009513173903, 0.0188701783862902, 
    -0.155525910627485, 0.386234388178982, 0.386359231366217, 
    0.282073398603928, -0.380636984078365, 0.409563901710436, 
    0.521417053575807, 0.0350718126352847, -0.264968329699441, 
    0.0635492635628908, 0.56237093570168, 0.0510916800010467, 
    -0.0119065808272523, -0.0163863315980258, 0.45750860145398, 
    0.0957751970664313, -0.0181020867194997, 0.152060344847646, 
    0.422846612709204, -0.0293795340812764,
  0.44031137175615, 0.073733960723986, -0.0386522208554298, 
    0.00263262731068524, 0.381203693365487, -0.00445449111246644, 
    -0.126578585328496, -0.143810821951275, 0.447212166927477, 
    0.226217154297848, 0.0230185976486418, 0.222003584614903, 
    0.312868704471551, 0.139674794711539, 0.0557591051805992, 
    -0.0618305387440826, 0.149077949405412, 0.293567110733116, 
    0.137579068056485, 0.0629121658272581, 0.0677498224172674, 
    -0.0493745447552974, 0.0712376409846261, 0.309828667232495, 
    0.295904943168629, 0.109300776337609, -0.0563959150107604, 
    8.19349500347788e-05, 0.224837549897854, 0.243048110208335, 
    0.145392013514028, 0.068595602420897, -0.0265983565005434, 
    -0.0104669177153945, 0.0344170446234954, -0.0123779392347117, 
    0.0276847822852146, 0.00403702061615482, -0.0603915791078099, 
    -0.0611749539421196, -0.188300636647891, -0.109992934427857, 
    0.017472543639594, -0.0736462780259685, 0.0455291805427894, 
    -0.0921980622396866, -0.0141928241480685, -0.0498607273237613, 
    0.0402752452218052, -0.175789122443538, 0.0901042289751839, 
    -0.010943235491593, 0.101425534895325, 0.281497523914889, 
    0.155702440048385, 0.0551223824235062, -0.0978775299694246, 
    0.0950702626712082, 0.292475391493703, 0.224018533220403, 
    0.164140019513955, 0.0482463506264205, 0.368644827608944, 
    0.469692403624735, 0.194650458016881, 0.0106484224702613, 
    0.148238948451215, 0.279269883144636, 0.301826024274668, 
    0.697678199140872, 0.674698046155872, 0.194408620781438, 
    -0.274652800440483, 0.375937640793237, 0.664408308947316, 
    0.0900614444485285, -0.00107037960686589, -0.199746709163002, 
    0.510140650150938, 0.364069799436129, 0.0691350122541322, 
    0.0323363955745076, -0.216116219156057, 0.430378614550191, 
    0.238963680708425, 0.110322861966124, 0.201522577261711, 
    0.237100784123033, -0.0112529707002835, 0.618445906015784, 
    0.194040696290732, -0.0301841087505517, -0.0343210224435577, 
    -0.034223822928589, 0.0617538955856453, -0.0614520112335931, 
    0.0421017633865701, 0.0869619865219281, -0.071454587861196, 
    -0.0431877777609625, -0.0395141193821177, 0.0171340981460007, 
    -0.0418245372027115, -0.00487368681034632, -0.0214043317175992, 
    -0.0154200859642058, -0.00609183106711664, -0.0117737672092373, 
    0.000276037327215956, 0.00332171954585124, 0.0761421539056693, 
    0.137016936925104, -0.0603768745708208, 0.290151786665913, 
    0.348509677647733, -0.0396451327337461, -0.256081632219112, 
    0.135956902961237, 0.569774234651261, -0.275452922896807, 
    0.32835094586778, 0.783951292500739, 0.0653173063391734, 
    -0.109977352377743, 0.0330862253033263, -0.0456024727500254, 
    0.614865051550572, 1.13297754361023, 0.426188629775906, 
    0.0220997360956916, 0.313254172498235, 0.381078828382854, 
    0.0788744777831853, 0.0435086978828588, -0.0738470755594494, 
    0.095105403270866, 0.16687588762746, 0.109080122173328, 
    0.0864566096894867, 0.0698025846372363, -0.0188899690173565, 
    0.0865990962128745, 0.119197981995811, 0.16640673634, 0.244761133240734, 
    0.0859023795510927, -0.0134055853266159, -0.0499554806199443, 
    0.298944306595935, 0.0714820962465371, -0.0311308098211151, 
    0.1854339017003, 0.196005747687132, -0.185341320945112, 0.50877861712012, 
    0.644826958138409, 0.154465713583128, -0.17628504336075, 
    0.293384786162871, 0.399347167078031, 0.13916454187316, 
    0.0892275156848066, 0.0471731309724104, 0.072439830407206, 
    0.0423404151360048, 0.0426111991161569, 0.061508285601628, 
    0.0795185797462894, 0.0985782701624561, 0.0315030062440414, 
    0.130651866100984, 0.115701263849293, 0.0349951860288786, 
    0.300331945274477, 0.267486499599367, 0.0786228507249306, 
    0.0604172496869778, 0.266179630940094, 0.140282343903334, 
    0.289468180712068, 0.493717373224583, 0.197471780307481, 
    0.085547416812836, -0.317840987295267, 0.00965208588459322, 
    0.568276577367328, 0.136430192582535, 0.0698348627986708, 
    -0.162268322373214, 0.463325546308894, 0.24211583231206, 
    0.0612102619069174, -0.13690421058135, 0.0860292507834704, 
    0.239939226030183, -0.0118397120584711, -0.201506836245658, 
    0.358403639612294, 0.230673411950174, 0.0653566489704549, 
    -0.085389836726583, 0.0736964214827046, -0.0995587619480975, 
    0.0497230804756081, -0.161330196038753, 0.0246407510331147, 
    -0.180801006650973, -0.024075731661475, -0.0897620823662738, 
    0.0410813288471164, -0.0421249688076549, 0.0359096319766541, 
    0.229210372342321, 0.103303199543992, 0.357347587208985, 
    0.330946557328748, -0.144780909660413, 0.37125448886483, 
    0.237216724742409, -0.199807827541844, -0.032506788981191, 
    0.874944674347365, 0.0700853469329471, 0.0267956786337618, 
    -0.0690386637050438, 0.573915360508243, 0.0692466974732229, 
    0.249901646718775, 1.10807341588328, 0.152733712376366, 
    -0.115068823842951, -0.113453930433394, 0.0892531559421778, 
    -0.0921434462178892, -0.0917935212773495, 0.0465259121807902, 
    -0.0044939415520949, -0.032045006632989, -0.211667850521188, 
    0.0713430494749417, -0.110219541206833, 0.125881333285607, 
    -0.235738502721031, 0.0425269748377803, -0.211003073467812, 
    -0.0298144193930593, -0.160761312698763, 0.000114154339692391, 
    -0.189477226110422, -0.0231417475790088, -0.053946865723827, 
    0.00318429384397297, -0.0546428050597529, 0.0169889501682588, 
    -0.0492034389949474, 0.030787658745397, -0.12080105271984, 
    -0.0185332153111706, -0.104791554074637, -0.121891073032908, 
    0.055550268386617, -0.0173178620583299, 0.0159494668866328, 
    0.0166815807526639, 0.0217711510034556, 0.0161750640261411, 
    0.0452704121295218, -0.0427462855159375, 0.0178608217122014, 
    -0.020894001336251, -0.000423435135030972, 0.0311471907404905, 
    0.0171057899424727, 0.00129104844366565, 0.0539228625806239, 
    0.0814967375530279, -0.0256724870661564, -0.0442091696269276, 
    0.210579750903221, 0.0745854209600687, 0.0958264140154012, 
    -0.163341667975126, 0.657388529840276, 0.22172383402272, 
    0.106031392493806, 0.600609939139273, -0.27242147663031, 
    0.336585421562903, 1.05788405027696, -0.0164753554336897, 
    -0.12189633178175, -0.0109992708933919, -0.12697145438388, 
    -0.0317655964758728, 0.0618283789995372, -0.130889152361087, 
    -0.129515058264868, -0.0407990234964838, 0.038254309088351, 
    0.085899323432848, -0.152291737985246, 0.172454208121642, 
    -0.367559339814671, -0.0269494392115376, -0.157305553891271, 
    0.0551317844507061, -0.372916896012726, 0.028984832488172, 
    -0.53230556810314, -0.271549115287006, -0.0412155369674095, 
    -0.00500985350436085, -0.00574487043600962, -0.00430931307164598, 
    0.0157218531878645, -0.0172237475560449, -0.0201219998703992, 
    0.0131786267606063, 0.0630080776261602, -0.181005840113748, 
    0.216440688683237, 0.316352868536836, 0.1501456067701, 
    -0.089010569819953, 0.264867170534617, 0.273533018756705, 
    -0.00865344317907746, 0.421441582107779, 0.63794824388855, 
    0.112736127336467, -0.277172329124313, 0.388488187556602, 
    0.63596694652104, -0.300431589243682, 0.268938347802173, 
    0.988446794953187, 0.903127957704884, 0.474904581418972, 
    -0.0371395674252137, 0.709106252585139, 0.466676107120872, 
    0.102907373678643, -0.0320430436929378, -0.124636923152453, 
    -0.0907445119379792, 0.725093663372827, -0.015390359916944, 
    -0.0775732055393725, -0.0740083068078486, 0.525971215957129, 
    0.110371979235733, 0.0510928635646183, 0.0938565258287907, 
    -0.0568057986353363, 0.469208494789378, 0.172987590054685, 
    -0.0300013339302883, -0.0663898352895151, -0.197678550745914, 
    0.0171723311615694,
  -0.0895285657536853, -0.045816480464961, -0.0515807756931502, 
    -0.0663327647008615, -0.0326788965515297, -0.066983243396075, 
    -0.0349679274109705, -0.0149277884386244, 0.187556235681252, 
    -0.0964568976882726, 0.442395295703342, 0.153636184133331, 
    0.0596801304209158, -0.247919669485864, 0.160758236415305, 
    0.499541958005047, 0.219544762640228, 0.0477300069999822, 
    0.535454592412474, 0.155311445258037, -0.0109449011046072, 
    -0.402003760274315, 0.451306583347125, 0.61048000451653, 
    0.125453494535815, -0.118775393984038, -0.14949527182257, 
    0.605272503367539, 0.295972544193972, 0.179278792049084, 
    -0.239634652760301, 0.299820083104672, 0.294030769703506, 
    0.116764315982425, 0.048366660792074, -0.272812145028338, 
    -0.0505208960762573, 0.378723778610663, 0.218620242184844, 
    0.118117227071557, 0.168915356448494, 0.337117192484946, 
    -0.159764314754392, -0.089794778970374, -0.0852599626245574, 
    0.287474570490648, 0.0806254668872919, 0.14832158613397, 
    0.452426235865878, -0.105170184375094, -0.0902255962560119, 
    -0.123824568385808, -0.0171894588655433, -0.061992566884014, 
    -0.0551460674607437, -0.0774305637065041, -0.0806281193174592, 
    -0.0543163556044622, -0.0392061685575953, -0.0971424227219285, 
    0.0468263780716418, 0.0315571363924052, 0.0574745631899878, 
    0.0468027565131377, 0.0610712490391601, 0.0343145746557668, 
    0.0541208211393537, 0.0445182721826038, 0.0376667288009769, 
    -0.033971038587094, 0.297722454883465, 0.176095985878168, 
    0.0413819563109561, 0.0140236605641767, 0.177590195238264, 
    0.340122776471737, 0.384526823444568, 0.341869237696018, 
    0.0657632854577977, -0.298484157195037, -0.0162528646183907, 
    0.567521854841511, -0.0553747489397816, -0.234612494200313, 
    0.345268082024764, 0.356577991776191, -0.556438233637788, 
    0.428644165703617, 0.630487953610773, 0.0801527363250486, 
    -0.0788167212036006, -0.214699030712037, 0.0986919587891488, 
    -0.108472957467168, 0.0247728370381356, -0.166990211149247, 
    -0.0125320908309799, -0.0723402452485302, 0.0314618010722519, 
    -0.221293567391631, 0.0123547914101643, 0.106609071037482, 
    0.11864822285149, 0.143278250899096, 0.20138018033185, 0.295778272695709, 
    0.323548213653951, 0.203812897031433, 0.0494444311531373, 
    0.169013908555108, 0.527774975635082, 0.257197866774608, 
    0.040198535580988, -0.0760539214124367, 0.737269228743572, 
    0.268033391708375, -0.00678693032777733, 0.0115772361956709, 
    0.334324813731337, 0.320017929943502, 0.683368507985367, 
    0.456197709757815, -0.108574974458773, 0.158663386017545, 
    0.734978910901605, 0.615833914659133, 0.232068269570282, 
    -0.19676297417698, 0.345604587410065, 0.450351768923155, 
    -0.127393471503006, 0.0267269227596462, -0.260504187097035, 
    -0.00493082611695434, -0.308755063001815, -0.202488657694976, 
    -0.0172021970973363, -0.0950619265542895, 0.0590886261316057, 
    -0.230295095591319, -0.04788798944574, 0.0864865931875029, 
    0.24351421078258, 0.228495285885583, 0.171621401271774, 
    0.170350948919645, 0.179389364117177, 0.256173900880468, 
    0.336278820710372, 0.291148680139642, 0.228955215438297, 0.2016268106508, 
    0.185064405889253, 0.188019631079396, 0.195352146144314, 
    0.182965494441013, 0.23965302232288, 0.215178455464283, 
    -0.00713386596045984, 0.0570223019308334, 0.508753744643371, 
    0.337998725052155, 0.111145208330578, -0.137028019097145, 
    -0.203849477852203, 0.65337320061176, 0.387881482560037, 
    0.151901516404131, 0.148370999489679, 0.203617449619158, 
    -0.0747725872752974, 0.536594994280022, 0.0783043539409327, 
    -0.0106977550045972, 0.211361831752032, 0.0666798707364981, 
    -0.0227870127411324, 0.674458229558788, 0.120763288008214, 
    -0.0370800824763382, -0.147694351513393, -0.0571511752271306, 
    -0.124588813810891, -0.0816774600049083, -0.104000374436426, 
    -0.0788191729848934, -0.0926623986589, -0.06949666644747, 
    -0.026123067917547, -0.0964413645625678, 0.198099051998072, 
    0.00864525382590105, 0.129772412771797, 0.326499340588432, 
    0.13753243907589, 0.0257145668375141, 0.453576143527172, 
    0.130061326853587, -0.189993121975799, 0.301427249863298, 
    0.417530684033189, -0.176987556484742, 0.0188493888187864, 
    -0.361242907608827, -0.0623922616547259, 0.633176634680096, 
    0.735477557499659, 0.250402686659402, -0.0199520751024972, 
    -0.112265069983706, 0.371474468798169, 0.282240971938214, 
    0.0943654992444801, 0.0507274443109947, 0.0416631368981158, 
    0.042864845895986, 0.0521162856594286, 0.0670880007294768, 
    0.0556353900311615, -0.0182902088660376, 0.0338687057265786, 
    0.193389538617943, 0.200215894169747, 0.13013562069798, 
    0.0495585370965409, 0.0412582375616907, 0.452194840247566, 
    0.262953072438807, 0.0597126548331074, 0.0760464454061525, 
    0.264385208917225, -0.118515808986428, 0.560512196702639, 
    0.53080691528669, 0.138027279280623, -0.103883025165069, 
    0.427930157587935, 1.13912120253919, -0.10560658001414, 
    -0.338377127540715, -0.395941113657015, -0.0599956899571545, 
    -0.250903405305718, -0.162970708727223, -0.220281018741726, 
    -0.0152836284906254, -0.286841954189082, 0.029692576550244, 
    -0.206774718387841, 0.0109337554755019, -0.0298957095236253, 
    0.158741188562725, -0.0678109637202744, 0.0492170414146911, 
    0.0442085531792836, 0.0368840302453999, -0.256500691559312, 
    0.0179457918427339, -0.121466127471701, -0.17905013367972, 
    -0.0112760080292324, 0.025741716789043, 0.0123929420974978, 
    0.0297018734409498, 0.0670053727883847, 0.0440993130078468, 
    0.0209850488639841, 0.101536465545499, 0.0996422758398158, 
    0.0305597302222075, 0.00602766248871961, -0.0635850659737053, 
    0.572780911373219, 0.35779418892834, 0.197338172374506, 
    0.140080115103531, -0.281358500147261, 0.49393228652652, 
    0.37542897264437, 0.219872024293415, -0.234827502516616, 
    0.678931014146426, 0.328653353909531, 0.0309136226423491, 
    0.163588102452136, 0.841535506616729, -0.058671972879436, 
    -0.00487867785335319, -0.217320917958897, 0.560453457113733, 
    0.305173259601719, 0.0326696428932951, -0.233804957824855, 
    -0.0723015030252095, 0.439948272704917, 0.106335914395534, 
    0.0156159956919665, -0.175336221179083, -0.00488005229837921, 
    0.35232621467695, -0.128567308925913, -0.0762365661889665, 
    -0.0397023463947538, 0.178565533653382, 0.00212257903385724, 
    -0.12806399369111, 0.0468856759212398, 0.173431077024432, 
    0.0156788579077369, 0.0613231331364498, -0.072936042345415, 
    0.0570837518431672, -0.0618579340628156, 0.0190510908028924, 
    -0.0366692944099836, -0.01068143266621, -0.0127071438221373, 
    -0.0700307555644408, -0.0580372639692374, -0.0668427970527571, 
    -0.0261500580681588, -0.0391112349953578, 0.0696988956157075, 
    -0.0443940780061349, 0.0390556114239972, -0.0230638469441012, 
    0.00826110857496042, -0.0160806777367447, 0.021618329987468, 
    -0.0795262028597771, 0.0212767104450024, 0.0658819447966384, 
    0.0648925685612921, 0.144806317752789, 0.129927161391194, 
    0.0361303768685599, 0.177366683203338, 0.189016145102755, 
    -0.0598083717196796, 0.046883709584677, 0.443453555338231, 
    0.306054002838601, 0.36973681047726, 0.242264861517518, 
    -0.199813114379256, 0.670040097274169, 0.666140609296345, 
    0.350473270376719, 0.208394846614329, -0.123155020453887, 
    0.269794004403439, 0.724549503639343, 0.00688249370358215, 
    0.0591626919160901, 0.148249077007815, 0.600752781224416, 
    -0.0670976236739338, 0.355692040315589, 0.781338664138703, 
    -0.00868862547917412,
  0.717353947271983, 0.367815006267235, -0.138974856793473, 
    0.380601543576973, 0.488986662673874, -0.159021575108788, 
    -0.172041417800709, 0.0498587342377852, 0.448805158785904, 
    -0.0196670391971919, -0.106301111894357, -0.0634412711711966, 
    -0.186127374553637, -0.00443021766176557, 0.108037956848024, 
    -0.0741496416769873, -0.214319576440357, 0.0125569492313928, 
    0.010962464511997, 0.00435351616517194, -0.169427547415903, 
    0.156568075147119, -0.205430229886065, 0.0436203435473863, 
    -0.142663570300495, 0.0538243620364926, -0.258656816846645, 
    -0.0161495982530641, -0.337558731535957, -0.194700050555253, 
    -0.00403253012490429, 0.0260923690473041, 0.119709778440835, 
    0.108717919137173, 0.0734108022419547, 0.0831141145336393, 
    0.0589315181657438, 0.0612302233205537, 0.119157204110481, 
    0.0823391835363335, 0.133083050669857, 0.216042605147191, 
    0.226951673039433, 0.184078126613838, 0.168194748304434, 
    0.121005981968677, 0.133127953104254, 0.396009118651464, 
    0.261628878395456, -0.165286013476353, 0.447199865750503, 
    0.468393361830114, 0.318394409755066, 0.233702866761866, 
    -0.381006042883964, 0.162920635158925, 0.595047488350257, 
    0.0710564944254479, 0.289027188403472, 0.928204715636027, 
    0.0817800188373216, -0.00076070565488362, 0.0333229260785147, 
    0.0111956832274264, -0.0203968434715901, 0.0260603997059526, 
    0.00182347483337372, -0.312373960284278, -0.0632523352213685, 
    -0.133747236963944, 0.0314643422131111, -0.202761367512252, 
    0.164635330569602, -0.113711206383999, 0.103838853065599, 
    -0.222974851545463, -0.0037182316775637, -0.0791013200585772, 
    0.0758603045313882, -0.237547384213333, 0.0451739483327674, 
    0.0494132787233464, 0.050327338216903, 0.0724235431400318, 
    0.0769813331381439, 0.0517481848346045, 0.0610675346529291, 
    0.0728801433511113, 0.0571336411034107, 0.039294329762174, 
    0.182948995015467, 0.0888303556108688, 0.0609707579857689, 
    0.32960252361136, 0.218985743729226, 0.108195970968508, 
    0.490891100244999, 0.251648840227512, -0.147004550838614, 
    0.279389412726261, 0.495815658862086, 0.0851724993204117, 
    0.261143336057821, -0.216560795300904, 0.801231284528217, 
    0.13120452295377, -0.361437938086985, 0.33932492347843, 
    0.764404026859134, -0.283004127292528, -0.111669132945157, 
    -0.134517989114553, -0.0488525925778572, -0.0964404011310483, 
    -0.0586298869718651, -0.0707868901812131, -0.15017145880811, 
    -0.0377718677840754, -0.0840755899020739, -0.0926508746806401, 
    -0.0647167540708648, 0.0576783907452623, -0.16680450018936, 
    -0.0230141160093852, -0.148579660756388, -0.155711250939667, 
    0.0157805168497039, 0.0161928385608006, 0.123035789173362, 
    -0.0537925830264095, 0.101612268021725, -0.00397841093148947, 
    0.066708527138131, 0.104952527008475, 0.0106606232309006, 
    -0.0360690932167809, 0.05782262883851, -0.0144240577839368, 
    -0.117799932344812, -0.232882953769202, 0.195622429219901, 
    -0.296099408379843, 0.155597536033106, 0.682633227156607, 
    0.35884158091124, 0.459240889177649, 0.52824125006448, 0.530237460220701, 
    1.26200155221928, 0.413493373967402, -0.082228170935669, 
    -0.0115584039035722, 0.0518517237275237, -0.0368665632416497, 
    -0.0362050001638636, -0.0329143885862276, 0.086774959080545, 
    0.315567436824224, -0.0297704363892437, -0.104699518591797, 
    -0.130571772113918, -0.112127126712298, -0.106014631439133, 
    -0.127665703861354, -0.104914733755826, -0.117442076080097, 
    -0.0625211319793666, -0.103665839100197, 0.04026777490947, 
    -0.18382481617504, -0.0655754779105309, 0.341893014258109, 
    0.180040443549816, -0.105817508854489, -0.015527910811654, 
    0.41094883725536, 0.298942659431988, 0.119882121196259, 
    -0.00190225598920546, -0.0421530688595341, -0.156047722009493, 
    -0.00326658259936424, 0.104206337233677, 0.708446984233901, 
    0.427641653629348, 0.13555135717523, -0.330221415532413, 
    0.59978794245872, 0.212014471767322, -0.148952721837135, 
    -0.348698122112459, -0.0517368283420903, -0.150118499624842, 
    -0.250611331263192, 0.130069501146413, -0.208834603241153, 
    0.000636483003676802, -0.0440638021000426, 0.0626993649315054, 
    -0.237764587992169, 0.0427348118974262, 0.106631174466276, 
    0.117773538209801, 0.195694661699664, 0.229724504124157, 
    0.156531424484424, 0.120506026155869, 0.183408155196199, 
    0.206336271136615, 0.154373254047344, 0.132129873809705, 
    0.142653051691026, 0.162114776728888, 0.176560794070279, 
    0.175881874899146, 0.150505436105012, 0.151454289538611, 
    0.213487295275467, 0.200065299891351, 0.115437608057702, 
    0.0696441216201201, 0.172229366313042, 0.342939758643705, 
    0.258743279575847, 0.107020156650377, -0.0515025119825494, 
    0.400909970871121, 0.367048045635076, 0.189795739454515, 
    0.157777932565972, -0.269878524497082, 0.0959367702241696, 
    0.315552598082412, 0.252023663890255, 0.726900940823169, 
    0.464790920027238, -0.116398594544553, 0.493568687356157, 
    0.674365806376819, 0.244147689635153, 0.0517018744717297, 
    -0.105562668863275, 0.232299658938154, 0.737487538978481, 
    0.0712962969173575, -0.0573433201189577, -0.163584261936067, 
    0.0893504729284212, 0.374201235133905, -0.126158814956573, 
    -0.0935948112499848, -0.0807981375398109, -0.0840464441923858, 
    -0.0955795659751253, -0.0661528237340588, -0.0900650409014464, 
    -0.0690269557157414, -0.0449724202373275, -0.07772171674803, 
    0.0423727904966886, 0.141089836550871, -0.119707490905779, 
    0.175460240439119, 0.421238581512327, 0.190371477678391, 
    0.0520703984870488, -0.100219568205714, -0.0570561768513627, 
    0.217807661084938, 0.366159259388338, 0.193932218085642, 
    0.208944110457768, 0.471428481299727, 0.41829875679116, 
    0.768740967147592, 0.508982644771238, 0.191834042097621, 
    0.55729462566426, -0.109964303729414, -0.284408090151141, 
    -0.303067723306993, 0.0288139480507884, -0.332356321151666, 
    -0.0934055993054116, -0.27839412730907, -0.136436776306664, 
    -0.255249093073931, -0.144889535741583, -0.126128806323183, 
    -0.209504755072165, 0.0711434754159662, 0.0275400704171324, 
    0.091456716164362, 0.0963943337665822, 0.127608838102177, 
    0.0620803267331082, 0.0861835330497959, 0.106523524804303, 
    0.119087872712557, 0.0441589246738226, 0.0701110953697111, 
    0.095352355315817, 0.110313654549545, 0.123481496941828, 
    0.12690833849778, 0.102405359409025, 0.0985066244220724, 
    0.141894416012666, 0.119298553013629, 0.067730641508784, 
    0.176303534032718, 0.151824078834693, 0.0451762329579405, 
    0.302769499998739, 0.343757273115533, 0.172225288764657, 
    0.113020636019368, -0.149431646925065, 0.42344379859035, 
    0.365896861542056, 0.192335892485277, 0.203879892958987, 
    -0.15102201814885, 0.335941274735371, 0.900079013845389, 
    -0.106874907939027, -0.409850008135806, 0.0397939122447961, 
    0.606766485940209, 0.0451585055819991, -0.0875168640922836, 
    -0.0370599481370455, 0.0306254100526794, -0.0229946566996216, 
    0.0489517787307862, -0.0459190155495519, -0.00688797968918149, 
    0.0183472096828763, 0.038578438557204, -0.0780069961379078, 
    0.033257836578267, 0.139787721023287, 0.125034667678611, 
    0.135268816905857, 0.23602103360766, 0.237857956160517, 
    0.216307462908905, 0.24557999761681, 0.174398270290761, 
    0.0700603371619321, 0.376116013621552, 0.456949035981092, 
    0.195276077977096, 0.00382215550353272, 0.332635997334082, 
    0.394751260650867, 0.26716781696806, 0.401042865194283, 
    0.304360991640485, 0.09444209724809,
  -0.0172075831682148, 0.351692393296804, 0.362657700950859, 
    0.332002292832953, 0.427878467054056, 0.393632502422807, 
    0.231293767574752, 0.116890542278821, 0.329663000082602, 
    0.498506823786709, 0.308838545732599, 0.174186630771968, 
    0.0743425605575088, 0.093735443299514, 0.282449128442102, 
    0.158828151029709, -0.0130707959739584, 0.113921051982374, 
    0.30573480224388, 0.223364975949698, 0.16187564503398, 
    -0.192919107560549, 0.0330308583722278, 0.559148527537971, 
    0.141085164938712, 0.0046805797002733, -0.192292925140389, 
    -0.0470117632621997, 0.469781108587376, 0.481427708000995, 
    0.196970721763539, -0.016070967772437, 0.326143818452683, 
    0.148070030593038, -0.233294498015696, 0.672172310756638, 
    0.393266571989589, 0.328998598021961, 0.65408503287099, 
    0.130769119123415, -0.157661837898689, -0.0179824809736965, 
    -0.208457477181838, -0.0779100195111763, -0.0878315981812194, 
    -0.242546988388708, -0.0500310597000918, -0.072462741254097, 
    -0.189105580905203, 0.00598545057863106, 0.00675572943420943, 
    0.102167944264765, -0.0387222682523437, 0.0777504597102417, 
    -0.0730642437023238, 0.029318696657552, -0.139800533070148, 
    -0.0524977396765652, -0.0418594525856276, -0.139198432169984, 
    0.0592301768400217, 0.0152734081164634, 0.0534370814403137, 
    0.0371920228575854, 0.0416347331497837, 0.0140825194271775, 
    0.0243429740983216, 0.0400962265771676, 0.046307842037688, 
    -0.0152613640370849, 0.0695271208450775, 0.109041372333571, 
    0.103849155186962, 0.12944759497031, 0.180404632481634, 
    0.178970523328657, 0.161127545061733, 0.121416710846722, 
    0.0410326489726719, 0.318162912961155, 0.31797493100204, 
    -0.00883767048025573, 0.15022547964052, 0.536367145095585, 
    0.222456076294665, -0.0305902858729606, 0.443545666064699, 
    0.429467563229595, 0.193686124673132, 0.0855803899397725, 
    0.0121112321636946, 0.314617604400868, 0.602199133692413, 
    0.197481790517876, -0.337419303872638, 0.214168186349894, 
    0.435472451264859, 0.751605667999367, 0.366435173260006, 
    -0.232314008411985, -0.306760677703638, -0.0982739400504557, 
    -0.143775385463677, -0.177048031737008, -0.113432809593842, 
    -0.118720961719101, -0.139727274630651, -0.065418094772522, 
    -0.186634837436034, -0.0651517070164103, -0.0380135876581678, 
    0.0660302473421765, -0.0894443257666746, -0.0141232048072373, 
    0.0136034826205044, 0.031852375940855, -0.120863261855351, 
    0.0200251880298801, -0.0815143069929687, -0.129010559751042, 
    0.0530537880063014, 0.0198512625694605, 0.167835607566655, 
    0.129994500393788, 0.033856259457779, -0.0865520526861608, 
    0.00604744519968022, 0.139670046140876, 0.0911926567508383, 
    0.339673577834257, 0.437142194078541, -0.137037705849585, 
    0.323502041307173, 0.580287488582379, 0.40499320681465, 
    0.179741037451351, 0.0311222286280073, -0.448188685243385, 
    0.114915863560617, 0.734515208206743, 0.0171578561281366, 
    -0.0862150753820362, -0.0981727956956794, -0.0726705801808024, 
    -0.10147140006106, 0.0094408374158516, 0.0187963235356177, 
    -0.185000960100099, 0.0786520154731655, -0.135407379233215, 
    0.136152525445843, -0.0505327810462622, 0.106126946163313, 
    -0.165194554691477, -0.026105723546505, -0.0296502385064507, 
    0.058207965853926, -0.0420627063270575, 0.0889139455823846, 
    -0.287241466760546, -0.00581979189278575, -0.0450859419671332, 
    -0.0235633949955387, -0.0614276001610378, -0.00768012325647163, 
    -0.0528061680843583, -0.0518493189303065, -0.00977906923590108, 
    0.00344958643373453, -0.0730634850150639, 0.27018067539718, 
    0.0851971809265282, 0.000511210083176339, 0.0170743371070229, 
    -0.00327338192217383, 0.248868270356488, 0.309726625484738, 
    0.668970565753782, 0.265664221345856, -0.557687474391024, 
    0.0704632199320515, 0.850818162333222, 0.17185702585947, 
    0.125132179344588, -0.423302856441164, 0.229009631020323, 
    0.502563202281345, 0.420124779915568, 0.708153073034783, 
    0.404213942005842, -0.183718402007531, 0.171758152926323, 
    0.542463759344868, 0.165274678925427, 0.025173536089323, 
    -0.0476076395399234, -0.0334061114450956, 0.171389403337719, 
    0.102775922734567, 0.0209457516254528, 0.232754066512092, 
    0.225841729947794, 0.0654395023168141, -0.0641342501933808, 
    0.0928711633875111, 0.152277695040559, 0.00169597495263246, 
    -0.00912241044641948, 0.243819219088066, 0.119415564483072, 
    0.069458949318945, 0.112349207045517, 0.130541974922713, 
    0.0773033246831311, 0.138213543313337, 0.116731928483005, 
    0.0123010426928599, 0.19232078416407, 0.208258915462814, 
    0.0678244082747954, -0.00467906555761423, 0.0521887069359882, 
    0.00843726556390681, 0.0497295276785942, -0.0758035441230887, 
    0.0326638650052577, -0.0280223327053242, 0.0551539062691156, 
    0.067044891520246, -0.0563354619225685, -0.0874917395407312, 
    0.294913066090238, 0.205491216390804, 0.0785448211243796, 
    0.0755210126492376, -0.127215076301901, 0.539271074279673, 
    0.105201354687203, -0.159294329238252, 0.0592163491476343, 
    0.51032388541029, 0.192069164818315, 0.166965338111831, 
    -0.338868392570991, 0.132316051684276, 0.533537562980976, 
    0.280050454082401, 0.138715798319192, 0.182598617595384, 
    0.193679457311941, -0.16878979388778, 0.357756506649785, 
    0.555139096173179, 0.249683431741959, 0.0281718835874214, 
    -0.209403958667201, -0.126364661060031, 0.578955486658332, 
    -0.00723608557610064, -0.0743021621714666, -0.0523205103249251, 
    0.393228237628628, 0.147255655882892, -0.0134372746217476, 
    0.192827669696717, 0.367352644166513, 0.333361926661511, 
    0.147857592501507, 0.34072902098399, 0.612492296697035, 
    0.213766403146452, 0.0213481183989515, -0.160348451413222, 
    -0.00450084829438809, 0.328054290879536, -0.040058110550649, 
    -0.15109337954184, 0.0689658126626775, 0.225405689823516, 
    -0.217611264987316, -0.242896973062176, -0.106751241300591, 
    -0.213437831031807, -0.211630810426878, 0.126189424342485, 
    -0.219888863219404, 0.0408890081433762, -0.120376094928339, 
    0.0265244327175794, -0.257905319424709, -0.017357102165388, 
    0.0770482197993826, 0.0849765585399079, 0.128590535465385, 
    0.192752004109246, 0.177014630070439, 0.175483661360009, 
    0.208309613247849, 0.156154575282489, 0.170896124851729, 
    0.336261139884927, 0.192185868824412, 0.0867891280742808, 
    0.542039874234541, 0.368508103290654, 0.0584710004191066, 
    0.347482520597544, 0.491319865711218, 0.227664986198082, 
    0.303101374991982, 0.378276433781677, 0.100438214267609, 
    0.175768161641411, 0.653020634257267, 0.664214026836498, 
    0.249488269240494, 0.035726133488735, 0.293119399089653, 
    -0.286232739572479, -0.329757543221013, -0.299547872724942, 
    -0.154838121680768, -0.247293903973628, -0.264286498395023, 
    -0.0257491236226404, -0.288771428293376, 0.0674932281919449, 
    -0.256619632989011, 0.0888166183910521, -0.217360003946666, 
    0.0997561441698596, 0.129206797889581, 0.127321220755353, 
    -0.0797051693534354, 0.0406395336415292, 0.0600806835698831, 
    0.0655580594184583, -0.236832308417582, 0.0154522251005512, 
    0.0185254018269281, -0.214700595154045, 0.106584046510386, 
    -0.35992591688994, -0.0297441419818087, -0.284106317307425, 
    -0.119788694601763, -0.213152902744882, -0.141628948270069, 
    -0.0134280878841148, -0.386628722850414, 0.215378217677201, 
    0.441504098328671, 0.00514976528248273, 0.26251911360373, 
    -0.373509366301036, -0.102179942564219, 0.635419785653975, 
    0.311202922961382, -0.0415074047841221, -0.125313039145661,
  0.0530627235771317, -0.209364480124226, 0.00403020899531661, 
    -0.0824388751198177, 0.0396596378199867, -0.0168643222026921, 
    0.105684871384324, -0.181299369696562, 0.0550404128624783, 
    -0.231719341719043, -0.0663145528792738, -0.00120660983429437, 
    0.0604619430735515, 0.073532479462081, 0.0767534508300425, 
    0.0110342079687468, 0.117967343805194, 0.286866413655942, 
    -0.214057631755814, -0.0776641055245267, -0.30813120197233, 
    0.109512285675577, 0.569744759945203, 0.394643084469576, 
    0.0195976025097654, 0.621236406440439, 0.405217161605724, 
    0.136981200429673, -0.20661755220687, 0.222755479397749, 
    0.391993509377389, 0.346401626766787, 0.48518321979806, 
    0.196061639504127, -0.24616971077554, -0.00855880110767371, 
    0.523676970268224, 0.205196489063366, 0.096120422268924, 
    0.429163205583583, -0.100912261955675, -0.177483174703923, 
    -0.126660843075338, -0.103335409627423, -0.04947145409941, 
    -0.0166313656695684, -0.0278296750983402, -0.190592033513001, 
    -0.193245042614519, -0.099877877662269, -0.103188427133144, 
    -0.148477605088362, 0.0312180250583485, -0.023378739253484, 
    0.0785765601738719, -0.119448507264426, 0.0476026582344775, 
    -0.0620198603005383, 0.0556031261705776, -0.175276326888565, 
    -0.00618415787501793, 0.0945598452030571, 0.0270063215756993, 
    0.0527885751519144, 0.263048024228137, 0.128322037984543, 
    0.00592419666558328, 0.0304341346920051, -0.0425482708880296, 
    0.475696479860321, 0.296284032364323, -0.0382638165761992, 
    -0.0827197535744162, -0.291980530381713, 0.764173778951232, 
    0.417873402083074, -0.187728370938347, 0.617683042223525, 
    0.678599954859489, 0.133342514548818, 0.0805261590027658, 
    0.368388446590686, -0.306000228047106, 0.235263658469364, 
    0.615254575086618, 0.379575447958438, -0.13706822362431, 
    0.992227019137241, 0.255791672325642, -0.00944959534866086, 
    -0.329258050271962, 0.0420422079600841, -0.41795251667048, 
    -0.140335441151828, -0.281563252436881, -0.269652970192657, 
    -0.112233251442523, -0.293335825644266, -0.0965104321451952, 
    -0.225608922467112, 0.0283438966030871, 0.0644413683874864, 
    0.0557824670769925, 0.0556873159061668, 0.0855413641555903, 
    0.0867530075015515, 0.0818119439228764, 0.0633235921658747, 
    0.0298986373141214, -0.080941937912635, -0.00510881724394553, 
    -0.0799884459168851, 0.363901234078657, 0.557420326094942, 
    0.338716682400656, 0.180389997271045, -0.376308800642657, 
    0.263347189561875, 0.411571872237395, 0.0385546319705174, 
    -0.0311001164291787, 0.477425174177332, 0.724290090697404, 
    0.362625252337825, 0.070867808200292, 0.208120995238677, 
    0.592401360757686, -0.0701803757976167, 0.639276369654607, 
    -0.00519068233492517, -0.328760759116788, -0.227436017181975, 
    -0.062275510916891, -0.240254522784946, -0.0462713278398876, 
    -0.220641232157869, -0.0459591661451195, -0.227504657717346, 
    0.0107084412268262, -0.193681408126921, 0.0593508084008727, 
    0.0899010600973264, 0.086522991055682, 0.124826862652642, 
    0.167468047515298, 0.183868078660868, 0.150851371140849, 
    0.081105866448295, -0.00867457204757738, 0.174478088295534, 
    0.417469598029592, 0.152698311321062, -0.00258395569033125, 
    -0.135897444320164, 0.273569810035075, 0.471480770863316, 
    0.112115184167548, 0.187259343007468, 0.771038271300344, 
    0.482957945467583, 0.289204336129461, 0.167160476469491, 
    -0.155196020398276, 0.0263090441583077, 0.207652435342737, 
    0.0390221665346029, -0.0581418717777228, 0.118692099770924, 
    0.244805829858559, -0.126388577433017, 0.0198341223215313, 
    -0.356710784449967, 0.07936220638385, -0.111507618837121, 
    0.097853652387577, -0.146129466657064, 0.142879540022568, 
    -0.26369356587233, 0.0407848747358154, -0.409069088790997, 
    -0.12801156936352, 0.0193883320229338, 0.0793825853156806, 
    0.0574718688783557, 0.0480743261945538, 0.0543167518089931, 
    0.233843822567416, 0.17785666419172, -0.181962678037139, 
    0.243565327182247, 0.548778723604561, 0.0611688206239951, 
    -0.404963555434353, 0.389273277795396, 0.729492645532508, 
    0.361308118973112, 0.21426366439778, -0.236007692678476, 
    0.592426518626866, 0.404852514685158, 0.532491644658046, 
    0.520059048314963, -0.318725732207227, 0.504382863601492, 
    0.44082422264016, 0.0577837518343185, -0.0765566029354777, 
    -0.0750304355542159, 0.457373588619594, 0.364317053945539, 
    0.111246109326933, 0.150261769657863, 0.218661079935199, 
    0.13596166687163, 0.0595504321013221, 0.0546701780287723, 
    0.184930161683524, 0.161800223992595, 0.0377895074070812, 
    0.136281303821257, 0.292600400582123, -0.040393849399469, 
    -0.175706218674941, 0.368517437438774, 0.399476744300962, 
    0.345174874221005, 0.0954867269600521, -0.171297645933329, 
    -0.222087570603357, 0.216415641521985, 0.522927623935103, 
    0.187454288109376, -0.182680901599917, 0.153982108579573, 
    0.531155093280886, 0.13244039454135, -0.134155091774331, 
    0.200189675446409, 0.371192358165165, 0.0401031086595069, 
    -0.161939242556657, 0.147636315452468, -0.0977901125500989, 
    0.0674832157252635, -0.117593152052781, 0.0311741552005454, 
    -0.310010441834207, -0.0696211290201688, -0.176493046939905, 
    -0.23182256695347, 0.0242796538448386, 0.0935097296802508, 
    0.132956296152128, 0.134866715512524, 0.274198446508283, 
    0.375826849294712, 0.21053281065895, 0.0353169847933448, 
    0.131907242740655, 0.398476855687958, 0.330774972368612, 
    0.219752087217855, 0.182978182656167, 0.188004364382042, 
    0.196270109128545, 0.169268756572693, 0.159558238541286, 
    0.205146689119698, 0.213989049018146, 0.177669762694749, 
    0.180781787596409, 0.187356653776691, 0.139540197596394, 
    0.106575470789493, 0.142216308246223, 0.275306702944194, 
    0.38560934055443, 0.148756920998966, -0.155743941535725, 
    0.0995420965902015, 0.425481200519074, 0.0762029910804811, 
    0.304780652683844, 0.567362436669911, 0.141165092998094, 
    0.278656591408128, 0.784066593646621, 0.127125642308232, 
    -0.0686000987201573, 0.243941232618117, 0.35524785005235, 
    0.0514005574608784, 0.0261124348581947, -0.116514427907484, 
    -0.242190030941978, 0.219530010099971, 0.217556300700625, 
    0.324029048778325, 0.269607620517735, -0.140228013213566, 
    -0.226664963244363, -0.104322463002906, -0.19498212584295, 
    -0.138982030717692, -0.195682534759356, -0.133674764916173, 
    -0.12832119384953, -0.181675086675376, -0.00687342967691096, 
    -0.185477855719496, 0.0818412176868082, -0.1161082996316, 
    0.00877307986414196, -0.0346461448958089, 0.0383774260592526, 
    -0.0510329646510185, 0.0763470692969403, -0.142177599455991, 
    0.0496549225657599, -0.112366185874528, 0.0677601080902736, 
    -0.0257691356962467, 0.113076424738771, 0.198444659772002, 
    0.105985084903702, 0.0397161251158693, -0.0168228765445775, 
    0.0589309436269873, -0.028328360505719, 0.343002963689558, 
    0.383349758775937, 0.114052124120124, 0.0867706891858816, 
    0.692470639413546, 0.153589915741624, 0.0767426237232347, 
    0.169066999213901, 0.142977010479195, -0.0833586735019622, 
    0.86239536786698, 0.184353224506156, -0.0657602903655638, 
    -0.0999346945647863, 0.512562392587948, 0.377025656115251, 
    -0.0320994009999845, -0.315245588276609, 0.00848072754284332, 
    0.371248499788321, -0.214640792378317, -0.214416829320086, 
    0.0655075812771121, -0.261104338008173, -0.0277818029340669, 
    -0.18913980298588, -0.104234910720393, -0.180437835344051, 
    -0.119203060407494, -0.0400003314649066, -0.16330847449822,
  0.323009559101788, 0.326539100201868, 0.0880784601327958, 
    0.170482797586274, 0.409414799945852, 0.184658173996464, 
    -0.0665658388233411, 0.325737918278802, 0.197203068160403, 
    -0.0332828324379723, -0.148274946470854, -0.0182928662852889, 
    -0.123168333821857, -0.0503236562176876, -0.123644456986277, 
    -0.0815516933439828, -0.0362902508328418, -0.10477547775781, 
    -0.0197200108553668, 0.0830903824477989, -0.146855732159561, 
    0.143479166780978, 0.275869580637587, 0.0567357743840011, 
    0.0171961940615905, 0.0423245361188141, 0.22048171592624, 
    0.699920994957793, 0.00737739577565108, -0.231186873281736, 
    -0.0850342501429891, 0.0914945440110273, 0.657841977828196, 
    0.605211503757616, 0.102151285444638, 0.550465510951075, 
    0.661475057702931, 0.311524032294442, 0.320306922071327, 
    0.664402010658349, -0.0650111873212491, -0.130274755308142, 
    -0.00183456633508758, -0.181569949902698, 0.131981903165473, 
    -0.168986520636504, -0.00119848108244043, -0.0554097241666139, 
    -0.0594095972729917, -0.0191357424223956, -0.22646637666766, 
    0.0847973628731514, -0.165795392140093, 0.0194426317755842, 
    -0.0514433623656879, 0.0783485756901977, -0.204623120046149, 
    -0.00504601280735908, -0.230298097362644, -0.182755040782677, 
    0.0461382268751142, -0.121132560362343, -0.0484476534367866, 
    -0.0192185796288989, -0.00865758788458887, -0.111011024345362, 
    -0.00947034164111234, -0.0292507178143028, 0.0378651767636401, 
    -0.099113029748871, 0.0334645761663154, 0.0579216478060378, 
    0.0554246571910135, 0.0607060274127486, 0.0694270295612148, 
    0.0580630297526007, 0.0549740464339909, 0.0844918842912958, 
    0.0672101154874612, 0.0096928071453445, 0.111575687500858, 
    0.144959860055769, 0.103583367407302, 0.22097552754273, 
    0.284552149783537, 0.126467673028308, 0.134283436149044, 
    0.402794994007502, 0.207673248397139, 0.050654537275506, 
    -0.0914738755784066, -0.177970547711229, 0.438687876730472, 
    0.452842452193016, 0.262594069150147, 0.260278465458857, 
    -0.274214250135832, 0.639196606549317, 0.234447006644978, 
    -0.0195848580571578, -0.0703709825454677, 0.60779150809844, 
    0.223414062718175, -0.144289729429686, 0.199474900426253, 
    0.403362475755965, 0.610898685798744, 0.157973713598958, 
    -0.282363887300492, -0.254419544922008, 0.119459009101858, 
    -0.282455403670866, 0.106303644498975, -0.27204893790929, 
    0.0951894693632412, -0.241320563187764, 0.0892475520663119, 
    -0.208072724746356, 0.069959619517885, -0.272449063370653, 
    -0.0286400087219952, 0.107284847948398, 0.141606809114984, 
    0.0531555220615708, 0.215442017736091, 0.410622237916707, 
    0.21160876405192, 0.043711920690843, -0.0499163252361613, 
    0.483115479863328, 0.339426070423302, -0.0598358571395485, 
    0.278072520199824, 0.641272055398034, 0.141540560299556, 
    -0.11000965989984, -0.0277034591380496, 0.512531139137048, 
    0.440055129699898, 0.232282907569051, 0.098244056751461, 
    0.0480372194131925, 0.187734214179706, 0.516404079808241, 
    0.357880022410839, 0.102703644992386, 0.0273371565220672, 
    0.511964321171155, 0.360393817268777, 0.0421709778809815, 
    -0.120121563086401, -0.0714413977706349, 0.535898047631615, 
    0.153482540130959, 0.0470154924385719, -0.121151295775281, 
    0.0739525082583129, 0.335578032534498, 0.416213107886948, 
    0.227333734567368, -0.00803285726215677, 0.528153567280364, 
    0.366248356655353, 0.162649435149038, 0.11512768415071, 
    -0.306065029512489, 0.243195047951173, 0.869296352235591, 
    -0.0842868441227027, -0.122659354245014, -0.154337917149773, 
    -0.194413926535226, -0.126544247068429, -0.158448966866041, 
    -0.144211926699693, -0.0883267760669729, -0.222565213772874, 
    -0.036565011478482, -0.261231068863905, -0.0796280876665716, 
    -0.0221216623758692, 0.0174075775682723, 0.0999257452712846, 
    0.0965770822485678, 0.00819702617934821, 0.0824591736278744, 
    -0.177201259276885, -0.0180536193696338, -0.0418528613316299, 
    -0.0711894568422971, -0.00509077517878327, 0.0495939953927247, 
    0.0566575199198171, 0.0644863484776725, 0.0839098361359047, 
    0.0572843488323279, 0.00865957749580719, 0.200869325414682, 
    0.0866440679002078, -0.193069860160467, 0.0979912170006413, 
    0.40402089159009, -0.0182977912367414, 0.171769962532485, 
    0.593844943279635, 0.294115449806399, 0.0810989054072471, 
    -0.135291758160844, -0.260436302381582, 0.385725362387171, 
    0.429034169414382, 0.139079041197462, 0.0876507621104484, 
    -0.297905088250856, 0.0679869820595554, 0.390437643384671, 
    0.666239316480086, -0.0431541999499498, -0.429634249693347, 
    -0.172178440752612, -0.137857417319865, -0.359683309422193, 
    0.0943963802236566, -0.303820005239653, 0.133806967921644, 
    -0.373796789879202, -0.0140584282857482, -0.337068041696548, 
    -0.273389503322995, 0.116033880275477, -0.164628096707999, 
    0.165307484192267, -0.0746873783894522, 0.0481995394129611, 
    0.218583502026711, -0.000899766532621402, 0.134598283757896, 
    -0.0657774344454226, 0.0188468212969951, 0.0324582762735746, 
    0.093041301431955, -0.0188742972535945, 0.0276200356450413, 
    -0.0553271820816916, 0.00702240787421449, -0.0451846603830482, 
    -0.0200758678572939, -0.00180587650440188, 0.0206070580306409, 
    0.0203881353308279, -0.100865616823629, 0.0407021224648429, 
    -0.103594442704994, 0.00129801003160492, -0.0940230258893591, 
    -0.00486574689948231, -0.086521692573314, -0.0129732521457393, 
    -0.0627351130898292, -0.0466285481322787, 0.0424893517317071, 
    0.0664317532087012, 0.156606962337303, 0.422135716326966, 
    0.128666509171022, 0.00762801144370533, 0.0158829899594704, 
    0.0772862087247047, 0.383176691764105, 0.160932911503382, 
    -0.467906939544151, 0.316889602589984, 0.501180856158839, 
    0.0294214393197724, 0.915267569390989, 0.617945185358765, 
    -0.219644978623435, 0.15328018943334, 0.966610953345215, 
    0.201906400287043, -0.0136248163942642, 0.0161682542049378, 
    -0.0126680465617975, -0.00461088290466036, 0.0326018706990293, 
    -0.00915399015905667, 0.0451767432532206, 0.0106628127371302, 
    0.0671610555659576, -0.0291431546107207, 0.140649118006779, 
    0.130850545891133, -0.0238732162188368, 0.199707129834366, 
    0.420048443549375, 0.156971908638292, -0.145897031464333, 
    0.298389173050649, 0.390556165304707, 0.0533018343415934, 
    0.12859709972295, -0.266884771124169, 0.384372489674248, 
    0.402494035248384, 0.32187500003828, 0.255775881540077, 
    -0.270478814970781, 0.417458179462457, 0.421380383923579, 
    0.0991286533407838, -0.158711392807843, 0.0727213066485669, 
    0.417955525485718, 0.14408820237137, 0.0861189155889311, 
    0.630019721951904, 0.192234635276829, -0.0488561134301962, 
    0.399459045116119, 0.22546804727182, -0.188895766557933, 
    -0.0187818549163446, -0.125669060825069, 0.0225193638664918, 
    -0.15388732134209, -0.0108273125149077, -0.0368589774173002, 
    -0.0468997816299524, -0.0570370265126504, -0.107357068835814, 
    -0.0943396972087854, 0.00933134916411883, -0.195267885739673, 
    -0.0716009561259307, 0.0248042492655346, -0.145954525213399, 
    0.0386556985266073, -0.0592118116469728, -0.0019190981364218, 
    -0.134172833008974, -0.0515178102490807, 0.116542617299224, 
    0.0675970257185668, 0.0318644572366466, 0.249373071299602, 
    0.125442573460984, -0.0386139448873167, 0.0887693968770705, 
    0.286189304707845, 0.135669056010855, 0.25000479405607, 
    -0.267021677320561, 0.317014005063154, 0.217550916734947, 
    0.211907033761487, 0.940651381292152, 0.534246496685009, 
    0.20075582068049, 0.145378701577035, -0.206766798007487,
  -0.274901442123229, -0.0483989252423462, -0.154743902667762, 
    -0.0479250013604733, -0.0941861401497644, -0.127494396573028, 
    -0.0784078085995491, -0.0994297743395811, -0.0972487528988496, 
    -0.128949155034087, 0.0659202898809143, -0.0589945623801604, 
    0.0621153217269561, -0.0341495169177468, 0.0348762059107973, 
    0.00601442273406223, 0.0859263639777227, -0.0316302754118772, 
    0.0775775131478806, -0.0842618646802795, 0.00352446577297034, 
    0.0511103073425608, 0.222936752170785, 0.0915251501188556, 
    0.0380650691608128, 0.0342998596069708, 0.146931054719625, 
    -0.00694379208234533, 0.227744818015635, 0.347108609456188, 
    0.264707140746406, 0.110973448796282, -0.538080485869028, 
    0.201816679541954, 0.59879876401005, -0.311026419388813, 
    -0.618503794126335, 0.259668243211102, 0.328886246310665, 
    -0.324473731161328, -0.0999483340496257, -0.120924783498854, 
    -0.0948597170565399, -0.0620919958555965, -0.111591410677694, 
    -0.0927819301183835, -0.100835410345945, -0.0352050599332766, 
    -0.134705858495603, -0.0217056936333542, -0.0300436245376775, 
    0.0593455519683828, 0.0902399403187953, 0.106933459567001, 
    0.0189038345744396, 0.0805056921758917, 0.0524949545286291, 
    0.0865639951032863, 0.0215520668363117, 0.0704391874696716, 
    -0.00310264000518944, 0.0317679569030025, -0.0149986201644642, 
    0.0214992840574664, -0.0409798042242772, 0.00852301499327954, 
    -0.00704077246610103, 0.0360765620770853, 0.0500995958720638, 
    -0.0336087645218667, 0.00861741960647083, 0.153797799034316, 
    0.107808239795896, 0.0307822974408264, 0.0944597619753927, 
    0.193904222639199, 0.231170567624627, 0.135297687029539, 
    -0.196790194025191, 0.0893555513588307, 0.446491227341845, 
    0.159758268554457, 0.0711814227626144, 0.129042841150279, 
    -0.0550392229820346, -0.477935019642389, 0.301862687035608, 
    0.802897794429542, 0.652904501083182, 0.0182952590575138, 
    -0.465684102462252, -0.253181524875152, -0.14108882471493, 
    -0.198268100135951, -0.074430199905598, -0.220206223001837, 
    0.0600370263010356, -0.140205401718464, 0.234266042824489, 
    -0.247285918647345, 0.100502199536021, -0.0363446257444697, 
    -0.0687303326819695, -0.287245740231043, -0.187535840275679, 
    0.01002430118793, 0.0812725360064894, -0.0877289246003447, 
    0.116622807273154, -0.327896124117781, -0.121819372881312, 
    0.0156918523875278, -0.0588755077802812, -0.0519724024791041, 
    0.0104482961136709, -0.0836355216488322, -0.0395487547873294, 
    -0.0243758935008481, -0.029490421672571, -0.048044662173225, 
    0.119837540642197, 0.106304815361696, 0.104175297969814, 
    0.00784669977737315, 0.32329714809541, 0.2581625776014, 
    0.113655673589878, 0.405456229318232, 0.24811791399574, 
    0.0262974648375132, 0.0914920004849147, -0.305220028954852, 
    -0.0890602916976514, 0.72149555383333, 0.203892434916256, 
    0.09500788867498, -0.33955162587546, 0.271457105860062, 
    0.604121566452049, 0.252067354692786, -0.0597910457928573, 
    0.329386621042712, 0.462732419704708, 0.217315348557108, 
    -0.0562600837058201, 0.364790225008286, 0.35532960994841, 
    0.0958726639610072, 0.00868277223312341, -0.144013486748257, 
    0.287959990521414, 0.290040494074926, 0.266232020389124, 
    0.199622986483589, -0.0658751811709628, 0.0745913504605709, 
    0.52432828764458, -0.0151128604722037, -0.121229068385993, 
    0.0486132147967228, 0.384569000474047, 0.00823083107570337, 
    -0.0694039416881154, -0.141278518961049, 0.365399901877533, 
    0.231049468432479, 0.301513330913032, 0.428531842018917, 
    -0.213216848962383, -0.173405225655851, -0.218532924879868, 
    -0.0638573186666006, -0.178592631912303, -0.142212375172904, 
    -0.0965921640435283, -0.151039696168708, -0.123566305704349, 
    -0.100231404269533, -0.154561980995667, -0.101587924985899, 
    -0.00966377149380914, -0.0186584844186266, -0.13346259223152, 
    -0.0130718257357769, 0.0435337180586741, -0.0869994052485366, 
    0.0508829524055006, 0.0227575472119829, 0.0619093082202813, 
    -0.0188055590459441, 0.0787555420552086, 0.0739880359550267, 
    0.0720584298018087, 0.0660302550974214, 0.0638737285880016, 
    0.0642243451222347, 0.0697361306951564, 0.0892532338398717, 
    0.0749326031953327, 0.0244400785659903, 0.0986371243136164, 
    0.11440809082739, 0.117621859258868, 0.290093785276439, 
    0.247159520179038, 0.0439420676410071, 0.237124818247011, 
    0.409055966795775, -0.119158473745772, -0.135513843669723, 
    -0.0751766892415512, 0.480513580496535, 0.0885429471280203, 
    0.0656987210230543, 0.73728288328847, 0.423614934894012, 
    0.052676445498667, -0.013744011959028, -0.389073118009653, 
    0.272440569004075, 0.381729777070454, 0.142987913180332, 
    0.0713068129199968, 0.198430504450135, 0.0282809124517742, 
    -0.058360363963685, 0.0776884496181435, 0.117782594608572, 
    -0.0591379804908286, -0.0462332038249885, -0.0454302057660018, 
    -0.164581935000043, 0.0286212750794169, -0.0820496990575103, 
    0.0170334482773197, -0.107917754922918, 0.0158773747992461, 
    -0.0158662869484146, 0.139063400919158, -0.150766333098571, 
    0.15341487463669, 0.254738501214606, 0.100292174346371, 
    0.00787569366828066, -0.033024358181774, 0.0231534088125838, 
    0.434582089288064, 0.0859467156854133, -0.0473127910161845, 
    -0.12198336806994, 0.406660131274718, -0.171465713750704, 
    0.342676515775927, 1.16084139144392, 0.621741621495563, 
    0.252545205977276, 0.271321063855041, -0.296173425889391, 
    0.954270618274609, 0.170660985661704, -0.00304746640377003, 
    -0.208052800065436, 0.245842681949223, 0.317880003772223, 
    0.461943778513375, 0.34900326324868, 0.134660451448974, 0.53173276616003, 
    0.212603357346629, -0.04153965061346, -0.157505408784001, 
    -0.00208057369316755, 0.274342270634674, -0.177637460923494, 
    0.051212127915927, -0.0942756425234671, 0.136053291371918, 
    0.0160814426598284, 0.233283850474751, 0.0714131547208161, 
    -0.0493739806039787, -1.45491442576778e-05, -0.0485684210640065, 
    0.152610070837355, 0.163634974806706, 0.108723110999218, 
    -0.0143296114083092, 0.19192853988913, 0.0736631178120048, 
    -0.118744975989612, -0.0262293588635972, -0.0385739235802834, 
    -0.0421848983124786, -0.0472267513421033, -0.0243603859833069, 
    -0.0483007427402963, -0.00415479781992947, -0.0462981930238197, 
    0.00555731740206253, 0.0514853113237869, -0.104686634697153, 
    0.254574369691897, 0.204333367165272, 0.00957862050466957, 
    -0.0274598589101819, 0.379519683983239, 0.245869975648075, 
    0.116871653898675, -0.16453470506472, 0.198473153856228, 
    0.416731229766797, 0.151039600002511, -0.0192673799305306, 
    0.335330959091892, 0.00416934809960456, -0.260378674436349, 
    -0.361039984763356, 0.0662929613973996, 0.328178272508894, 
    -0.120817779013386, -0.109044790900631, -0.079220121510084, 
    -0.112889838274184, -0.11331471173129, -0.0447093071363043, 
    -0.119113603887304, 0.00772828014740966, -0.0855296094940032, 
    0.064588472179966, -0.135294951842333, 0.0340624708961207, 
    0.105502171112308, 0.1153077924342, 0.15171877422074, 0.18017732218866, 
    0.144944566509607, 0.134060204489058, 0.190514001097207, 0.164479758396, 
    0.126086331882783, 0.208155835242118, 0.151579366480814, 
    0.257499034968692, 0.387849189421663, 0.154517288152579, 
    0.125867210107674, 0.625312406714219, 0.312020480739932, 
    0.0710813586551356, 0.278905481520053, 0.491885329990654, 
    -0.316416353948112, 0.197994945634073, 0.703466212830444, 
    0.468242929636772, 0.483746484422263, 0.352269008722257, 
    -0.0620554969317966, 0.471709866567651, 0.633542878439151,
  -0.0742478641219915, 0.138998206509398, -0.167046695404533, 
    0.104073772157315, -0.26234770814801, 0.00130742968725726, 
    -0.257612530034099, -0.14885558675776, -0.0297079263321961, 
    -0.216816226573878, 0.00466495609314305, 0.109966989871378, 
    0.130253147153155, 0.122859391412263, 0.138868439771329, 
    0.168277307811392, 0.215831563284737, 0.214058361508253, 
    0.155854528099327, 0.126463463678266, 0.141214921246612, 
    0.164955618935289, 0.178633827283079, 0.183415031398053, 
    0.19017476125928, 0.208393597835376, 0.240107419709115, 
    0.198289426647513, 0.0921985752581486, 0.205302208184622, 
    0.4414801631168, 0.16593397943957, -0.125341617227341, 0.110600990367652, 
    0.465961417437602, 0.212275048805084, 0.0635611810532125, 
    -0.0920596437008004, 0.00260984362994618, 0.579373825848937, 
    0.0303982026644842, 0.0178248463721972, -0.0239607348311404, 
    0.417735336579729, 0.101935089666252, -0.160481228225095, 
    0.712778714210453, 0.189192638908713, -0.216699876464335, 
    -0.248118752911659, -0.285740938387541, -0.311452242786979, 
    -0.00963982595687179, -0.0538059068716368, 0.102976900038676, 
    -0.317799966695635, 0.0279730719063548, -0.125456819717153, 
    0.076138828068617, -0.388530609229187, 0.00265884855247155, 
    0.0637946051344029, 0.12019571484492, 0.189204255768124, 
    0.140195343316463, 0.0620654264250413, 0.0877395653094017, 
    0.153502473088964, 0.137447340473969, 0.0678808734419017, 
    0.0799551493660373, 0.109161824213092, 0.11760877838473, 
    0.138264385709136, 0.16093854581322, 0.144151486567849, 0.14738381374866, 
    0.200142670661586, 0.165695784989173, 0.0816244960433282, 
    0.0994201328721134, 0.241575872109451, 0.297878463856681, 
    0.162145037591305, -0.0713492156758161, 0.252900676332917, 
    0.563774589253482, 0.0664772363756826, -0.13797554120652, 
    -0.0629456761118205, 0.574029709011905, 0.22241654800729, 
    0.107700430753474, -0.343949561061791, 0.127495857568638, 
    0.615767466504499, 0.0154415453489975, -0.168003431269665, 
    0.145276127774508, 0.560493627152885, -0.110480937569018, 
    0.053001610374134, -0.160645708939344, 0.0285315888923785, 
    0.0857604040004568, 0.359602565408121, 0.334137664094906, 
    -0.0591970306659451, -0.0912235974566303, -0.128092416567598, 
    0.221635513651711, -0.183878313128657, 0.130886285490711, 
    -0.125882598590197, 0.0716474238339396, -0.232215555614768, 
    0.0141481256851746, -0.145088894664907, 0.0238274713718638, 
    -0.376473789627957, -0.0328383836219522, 0.0461854891527408, 
    0.101706795594778, 0.131180175332359, 0.132940554902101, 
    0.0910787918880903, 0.0933755807879889, 0.155558157514617, 
    0.126710668708436, 0.0676192277145616, 0.13456290070735, 
    0.0837932428842054, 0.130430492639055, 0.358059901654461, 
    0.343633145403001, 0.151824408071438, -0.0666215986782685, 
    0.260898722265746, 0.463786733133689, 0.17897736265402, 
    -0.040429493405198, 0.455163250524978, 0.519191203781037, 
    0.196084255451552, -0.239980350342042, 0.510251227871385, 
    0.374103036160573, -0.0687717801491949, 0.261074275511069, 
    0.735463232205822, 0.0965266258444639, -0.323302945133227, 
    0.234321602384578, 0.5183707763878, 0.129613096223804, 
    0.0633121633045391, 0.0632866496258932, -0.156384109025398, 
    -0.108875953602499, 0.354666605679755, 0.462834817121756, 
    0.345569539677437, -0.0368930622525209, -0.245698408156087, 
    -0.359595688997942, -0.155728712137839, 0.188041075872299, 
    -0.0828222846799025, -0.168315683013622, 0.320289898707778, 
    0.0234513427941091, 0.171442321598754, -0.110488584790113, 
    0.144246211921679, -0.0890638423774357, 0.0833027819859041, 
    -0.375956289049713, -0.0454428988331997, -0.371125564633001, 
    -0.292326949372186, -0.000925223179204505, 0.0499128587933225, 
    0.119329803688372, 0.126729644810675, 0.111802220945795, 
    0.101598841252666, 0.0490157790247313, 0.0466167523237621, 
    0.124160086587804, 0.0675887960577276, 0.129315327736034, 
    0.161861673872079, 0.148122422519591, 0.157689924639188, 
    0.208744671032307, 0.209701216766806, 0.207042131738833, 
    0.251376836878418, 0.226586769438264, 0.200889967854275, 
    0.31098605259189, 0.244452829184373, 0.0353807800186194, 
    0.171408544976571, 0.57775657133759, 0.209345034640685, 
    -0.0471869222297075, 0.0659638851402289, 0.581577455515223, 
    0.130696937919652, 0.0611962848157974, -0.167345092778421, 
    0.452565139247399, 0.377182766617724, 0.263799113780021, 
    0.243788004516972, 0.0245035440460838, 0.760105862502623, 
    0.0814994633019359, -0.0283234281304707, -0.245575325582223, 
    0.429138626274518, 0.417677986290689, 0.183368101714824, 
    0.100041191349634, 0.412876101980685, -0.223773272595407, 
    0.452402971398669, 0.541902151219344, -0.163810781495096, 
    -0.196451269781259, -0.0537029540251248, -0.153666028149101, 
    -0.0650286242826305, -0.0204656255542426, -0.154250940560729, 
    0.0509931739878635, -0.0820587997752887, -0.162739537595518, 
    0.178662573235597, -0.0551354921191788, 0.173469516039592, 
    0.0140345021158481, 0.148017289315498, -0.155980689553545, 
    0.1371031180153, -0.250607477839822, 0.0155129431179177, 
    -0.24226435726994, -0.106802013127013, -0.0448266485548807, 
    0.00201692276105214, -0.0454080384103238, -0.00780065378668313, 
    -0.0479052016691099, -0.0150927119292886, -0.0868501330599619, 
    -0.0242091507066091, -0.096649082005097, -0.0659124301024742, 
    0.0139519647709241, 0.0650054404452399, 0.0482931305376627, 
    0.0577371114854449, 0.0453644813967635, 0.0410220343610974, 
    0.0681416699221774, 0.0670583170587184, 0.0483341658625659, 
    0.0666909129389942, 0.0677408280660029, 0.0763778991654806, 
    0.0738303018624902, 0.0741500069324253, 0.0785013190203302, 
    0.0780878644716805, 0.0848493326720527, 0.0984967776657046, 
    -0.0473891352793011, 0.0822604371648268, 0.408037588252139, 
    0.104782413507359, -0.0457086106721873, 0.42413556498308, 
    0.485483360046131, 0.241486845177039, 0.00449669485389197, 
    0.251954063413274, 0.440316763696886, 0.241795177590808, 
    -0.18396803444373, 0.877025690324926, 0.481017347305322, 
    0.0814614296221111, -0.391541871970193, 0.43490765233831, 
    0.670734413376814, 0.311434265818671, 0.158335661408141, 
    0.117078683898201, 0.0166940741210711, 0.352090229812627, 
    0.251583079890915, 0.0765114910951457, 0.021712578366398, 
    0.00275332245461063, -0.0198612760750947, 0.0339182767893027, 
    0.0536342329090965, -0.0692105322856322, 0.0285955802652186, 
    0.271443993794638, 0.246089094101927, 0.183447877834024, 
    0.142097143848068, 0.0456682711967846, -0.0987998001298847, 
    0.446031835972317, 0.237495841612285, 0.0528491128531536, 
    0.00395587212850479, 0.3565513587566, 0.197280768938302, 
    0.0281000584899272, 0.059602941778301, 0.340321072399162, 
    0.205573548428889, 0.0550840033646453, 0.26745615485123, 
    0.329475175644677, 0.144759818877116, 0.0907328950430482, 
    0.0939272423738035, 0.0983273569376867, 0.100133234726855, 
    0.0960838040784172, 0.10359062557317, 0.144917929178364, 
    0.126883265981595, -0.0875377291708548, 0.271053396673091, 
    0.265607491767087, 0.0450052378647906, 0.0291601446825438, 
    0.327282986190946, 0.347275120975323, 0.258139726034104, 
    0.129373561501054, 0.0936852452245293, 0.700852002339945, 
    0.200327048999815, -0.015708809190448, -0.234731232351016, 
    0.337423129216145, 0.666397062762894, 0.178810595160176, 
    -0.33619476776068, -0.0840810955808735, 0.555119343713661, 
    0.142572750670623,
  0.131935706824132, 0.050226261395845, 0.0324750165263093, 
    0.273082972313599, 0.23800500148193, 0.0773161027709175, 
    0.0157376134757316, 0.357233491864298, 0.285161333458248, 
    0.0718253748775695, -0.173212567222329, -0.0466022770332492, 
    0.472050846810503, 0.284449869611991, 0.0936314921623977, 
    -0.0188477142290542, -0.0943274645510158, 0.0772222661564539, 
    0.390429632803127, 0.461103337494485, 0.324951041494631, 
    0.175097132561968, 0.0599052297908137, 0.153204263153495, 
    0.160163790877446, 0.30571483004014, 0.660632018194534, 
    0.299399503994415, -0.0602896781318659, 0.141760962736277, 
    0.603012560697323, 0.178712325688158, 0.0986032680517017, 
    -0.192738986648458, 0.0965938632277693, 0.349510287158976, 
    0.0882612146903707, 0.234603554391211, 0.592235140087566, 
    0.242877863126084, 0.0316364008575337, -0.189237313177692, 
    0.0436875337592824, 0.290598887301396, -0.151613375332831, 
    -0.0865933151647374, -0.102995569454713, 0.394369018106133, 
    -0.176522891384563, -0.106645655140812, -0.27018428051649, 
    -0.191741559700243, 0.122872757408919, -0.164040712143442, 
    0.177530548711846, -0.134194144833415, 0.0436090412331637, 
    -0.0927943813936957, 0.0881920366245429, -0.332459596222002, 
    0.0107274409222887, 0.0625060513532637, 0.0571890384253193, 
    0.159354645155103, 0.225225277172469, 0.157869472547162, 
    0.115809555167781, 0.180391491781016, 0.189842645002528, 
    0.13823422343548, 0.179106056891829, 0.206605907880953, 
    0.208536321889594, 0.234738115083152, 0.226139592549099, 
    0.140922874378922, 0.18741728197137, 0.374443146628891, 
    0.224245003535669, 0.000450334237008663, 0.210183774251772, 
    0.525003535741798, 0.273653948144396, 0.165460684876235, 
    -0.2678679931035, 0.808251561023119, 0.181687944115271, 
    -0.267546589700985, -0.0761055581419348, -0.404779602262233, 
    0.322953612582472, 0.154000516888815, -0.10844212925012, 
    -0.118123094826436, -0.124103028238168, 0.112362829120876, 
    -0.0258024426356488, -0.179727021314859, 0.0876403040123035, 
    -0.00331087192597908, -0.197210433319413, -0.0204577240804505, 
    -0.618748298261821, -0.0963159777650679, -0.132332794965469, 
    -0.457516110184916, -0.00386123517390294, -0.0586361066207985, 
    0.0564257390157315, -0.459376244142953, 0.00160357069323623, 
    0.0110298159338934, -0.0519831390570746, 0.142178121100243, 
    0.057678418068291, -0.100130921322356, 0.0595708589739755, 
    0.305002823205967, -0.231362745465381, -0.0913675325545165, 
    -0.457401413367935, 0.59719991725218, 0.331488193917214, 
    0.0539780758061105, -0.0842329352213345, -0.257339296732543, 
    -0.0437865838307544, 0.651211550412255, 0.607271333672433, 
    0.114504797797259, -0.25646072653529, -0.025908258113446, 
    0.516933088257071, 0.241302249565792, 0.0734294039584562, 
    -0.0502476361349824, -0.222861208254609, 0.41287732807156, 
    0.480891636356957, 0.0552335458216263, -0.0236681506875578, 
    -0.370951368274302, 0.134099232289253, 0.319100811540022, 
    -0.0705762272837795, -0.158633771014171, -0.159938487932666, 
    0.268196471008808, 0.197042428055199, 0.0913808239460791, 
    -0.156791446643205, 0.131447234178813, 0.191206501629456, 
    0.232657483079725, 0.207537026438182, 0.0293905565198001, 
    0.394452418092722, 0.164068273840747, -0.013876719038917, 
    -0.00655052189548358, -0.251790398689574, -0.0104006215915954, 
    -0.164480623129169, 0.0415411008772374, -0.171257432079108, 
    -0.0101704038263077, -0.228397165512516, -0.149774283705995, 
    0.108662563599114, -0.228625052710931, 0.0284934810974861, 
    0.0781997312157355, 0.0828255629755866, 0.116539880612809, 
    0.139239443922716, 0.107199463036541, 0.107264191746835, 
    0.151870246051279, 0.119323891471069, 0.0662344915784424, 
    0.195678698595589, 0.179601959343738, 0.0464370052210071, 
    0.216442146491897, 0.421851238833112, 0.210703210785758, 
    0.0446391241056857, 0.133381676279289, 0.30190405075953, 
    0.208175574362597, 0.284321809354045, 0.323905908506141, 
    0.155338602326492, 0.618324615066083, 0.731543887772493, 
    0.440405371035339, 0.233188972264728, -0.566660351462555, 
    -0.0357109301995795, 0.465275737774085, 0.712483890427921, 
    0.414372307055427, 0.0209188068267962, 0.421212594817131, 
    0.267561518396434, 0.0645095479865013, 0.0497746533088375, 
    0.25783797407723, -0.239852223497592, 0.307305407558268, 
    0.217761459362181, -0.0126249661303207, -0.0515659544569024, 
    -0.0508156649697294, -0.0443960976678163, -0.0467870293031609, 
    -0.0483841744868093, -0.0317425153728845, 0.0418768739671576, 
    -0.167685878297909, 0.30128159988449, 0.214058319247519, 
    0.196789223076965, 0.183498400446034, -0.281465872043591, 
    0.316580631196084, 0.431723676060491, 0.107735945174879, 
    0.0223022355343607, 0.0512541754017828, -0.426416491812127, 
    0.563300347326097, 0.359393686033031, -0.020827711213519, 
    -0.0544587924188533, 0.410403549534375, 0.692607570091223, 
    0.354103555993408, 0.199691260272118, 0.555445415679902, 
    -0.0387288898577453, -0.176238470632527, -0.159976595722002, 
    -0.019773808226442, -0.116230136751524, -0.00276722536983774, 
    -0.127569333565109, -0.11730046778974, -0.0534376452671211, 
    -0.0540062827499749, 0.00123130306832527, 0.0151543826627283, 
    0.041682372892256, 0.0646152504038788, 0.0677527925198955, 
    0.0586299398784203, 0.0490769406347731, 0.061231336102023, 
    0.0569173619483757, 0.0309496699283725, 0.0667903933138037, 
    0.0438450818153703, 0.0574840236578399, 0.0562371610885381, 
    0.0652618792712242, 0.0286952595812361, 0.044487195784038, 
    0.0590722174989611, 0.0571451554811813, 0.0011876519477718, 
    0.0387779402886297, 0.0669713193591922, 0.222253057675194, 
    0.250165563698352, 0.122550938930492, -0.103754408872408, 
    0.239200563950798, 0.384829899605687, -0.0454522230062744, 
    -0.0215400370460949, -0.102440495457179, -0.112649337292946, 
    -0.0680355364411009, 0.848160284306564, 0.428232354127388, 
    0.00271833400121634, 0.595354194800539, 0.582314121577871, 
    -0.202407210563769, 0.778475095354699, 0.499702147690527, 
    -0.234720386510529, -0.222221316088107, -0.0114727381616324, 
    -0.115794681426362, 0.713629058058528, 0.457846785404121, 
    -0.0958688880189104, 0.693784372137528, 0.325500821258254, 
    -0.240551556168916, -0.0708211835409462, -0.123486346369551, 
    -0.0503811559298743, -0.17298041428537, -0.0747816683795149, 
    -0.0629335729417199, -0.0869148360293954, -0.118262710533187, 
    0.00171437304841515, -0.157042938711436, 0.0692399972740701, 
    0.151351769022499, 0.147117276845847, 0.447281180919766, 
    0.29146400591989, 0.049904170698818, -0.132148583618478, 
    -0.0389052079599559, 0.0926785461387582, 1.01436896110007, 
    0.0420853407665364, -0.305521154271943, -0.0527973422407403, 
    0.657100489941632, 0.467836304574449, 0.447913337997633, 
    -0.13589179658581, 0.536950009669775, 0.424024163969976, -0.170423849579, 
    -0.170612771003393, -0.130452432234158, 0.148747602151067, 
    0.0987377911660238, 0.188666244433745, 0.243665521946295, 
    0.047003571668583, 0.374779793081179, -0.0466078622505613, 
    -0.345382721393424, -0.154361157925528, -0.11246469576867, 
    -0.242365993548347, -0.0475389819104564, -0.187813093307082, 
    -0.0317086448107454, -0.260555161320801, -0.0858265412908102, 
    -0.118498364997496, -0.0505274502237836, 0.0488905155049935, 
    -0.0358416369914447, -0.00773700431893001, 0.0250753867735949, 
    -0.014248735131234, 0.0394211290654083, -0.0183578594291126, 
    0.0263170325866931, -0.00929842614906662,
  0.0105257004109294, 0.55075064653612, 0.36577215563069, 0.0989758610319381, 
    -0.158557723912159, 0.0653704886327937, 0.420129931644014, 
    0.285735967080392, 0.238228984136793, 0.176652157030426, 
    -0.209250708145968, 0.143627577632524, 0.44902286499175, 
    0.102741763842874, -0.189557653064766, 0.498494849298324, 
    0.473467317979228, 0.175775790977265, 0.0448451969387179, 
    0.369332768238251, 0.0371442760987804, -0.104338163232706, 
    -0.112924987967574, -0.0728312795512694, 0.0285288132843136, 
    -0.0289912162433496, -0.0440814277744855, 0.0183069810765381, 
    -0.0766982182070327, -0.0837682161280148, 0.0467611851815806, 
    -0.121932140799988, 0.105696374328145, -0.0939020642806514, 
    0.0698448101799894, -0.207041317224843, 0.0248081058839306, 
    -0.109099903471124, 0.0164614148662816, -0.216867554879924, 
    -0.0400873545950893, 0.0532305913636781, 0.0557716881668021, 
    0.0944937142262197, 0.139401566841868, 0.0950956044015604, 
    0.0602816999341751, 0.145301783993678, 0.152861497690655, 
    0.0945751082959243, 0.128909472260289, 0.096441976284864, 
    0.250654128827486, 0.126620375941262, 0.260797723763923, 
    0.714458253957461, 0.26216461668673, -0.186251892430295, 
    0.374213371947012, 0.527019589779947, 0.103580758673376, 
    0.0349071654887255, 0.0811735213730658, -0.10432312601144, 
    0.825630078858513, -0.0126825340323559, -0.13527595100996, 
    0.0708749273655961, 0.582014313529893, -0.10966674496826, 
    -0.199950314006351, -0.143554056145738, -0.0557834625691061, 
    -0.0701538987457934, -0.155591308505361, -0.211726966952772, 
    -0.191520209681824, -0.185801382705914, -0.213976128125972, 
    -0.138265269482194, -0.363130918706908, -0.193646686844071, 
    0.200504903082284, -0.29166444066774, -0.0321348656998267, 
    0.0974953459315507, 0.0733446667749216, -0.0569948990377149, 
    0.0671502388023117, -0.355785206807238, -0.0569541599712446, 
    -0.0537327934123742, -0.0433912955304346, -0.0387770504481981, 
    -0.0453573763033769, -0.0439472583494848, -0.0568032235749675, 
    0.0485582745781437, 0.11131844677153, -0.229031861447171, 
    0.334627604107884, 0.127791837342729, -0.0329946076743541, 
    0.078562330094224, -0.201683849097204, -0.0517527677168175, 
    0.771279124814228, 0.414679000225131, 0.348383130475682, 
    0.743819895525364, 0.215712224228214, 0.040494632297697, 
    0.023204125055518, 0.0427877629640892, 0.0415869328540788, 
    -0.0359334573117254, 0.0498410071739466, 0.0708620499070888, 
    -0.00866491435590565, -0.0304716784434252, -0.0367420488333272, 
    -0.128700452029492, -0.000790543563681592, -0.0545707828763557, 
    0.0083575624388135, -0.0228880526214374, 0.0460665836235955, 
    -0.0903979776390813, 0.0310391228382133, -0.154938201559502, 
    -0.042223965982722, -0.0166692010690704, -0.0319072813295358, 
    -0.00936836208492731, -0.0227618871306267, -0.0699223092727655, 
    -0.125320332011208, -0.11111122644177, -0.134629042719401, 
    -0.132108528218522, 0.125589745575649, 0.314160943124233, 
    0.368385447066147, 0.061186114399414, -0.564366684708631, 
    0.899574439662757, 0.455204444174545, -0.0187777256846305, 
    0.882011395192919, 0.618304657905809, 0.151840848772759, 
    0.102732749315119, 0.0225339732899333, 0.067654564746186, 
    -0.00725506048871483, 0.0227266963959057, 0.0168514597176707, 
    -0.00124541687385768, 0.0734717838824649, -0.00701076884690768, 
    0.0742400903798377, 0.00961715603676416, 0.0375998174629791, 
    0.0615877673436266, 0.0556564143857762, -0.0221829430065232, 
    0.0354629589131166, 0.0195183502355642, -0.0159950364015753, 
    0.035454266000533, 0.0474008083902944, 0.0619931635443827, 
    0.0157206012565125, 0.0505940265453615, 0.0401210541959529, 
    0.0515624102526384, -0.0153250946969782, 0.032425427362187, 
    0.00605350374382491, -0.0211399633044613, 0.0491750098076218, 
    0.0724730741002433, 0.0670925823918338, 0.0742847349338657, 
    0.12177911140983, 0.0981816890671285, -0.0925488341049986, 
    0.171322874120827, 0.25265131411724, -0.026173526394829, 
    0.166940949355926, -0.0907043063597013, 0.619805448566216, 
    0.630539075463964, -0.0347172545412156, -0.0463742598061732, 
    -0.300469690605125, -0.131213447101496, 0.515580097440182, 
    0.590260172374334, 0.181932622224681, -0.0360783410519704, 
    0.052509651400885, -0.24925565307008, 0.379266738636636, 
    0.0661780530313874, -0.142371073269795, 0.605870992288372, 
    0.374047787449229, 0.0964430038205771, -0.0491210445806468, 
    -0.177235510518004, 0.185098780468255, -0.0908879852697241, 
    0.0774412744670338, -0.0887684219353312, 0.0991055402417201, 
    -0.251607965690948, 0.0602061338129049, -0.312070850382751, 
    -0.0602651880680149, 0.0445931214581349, 0.158122060161249, 
    0.193796251498583, 0.21765904743586, 0.271816359559099, 
    0.230663500411876, 0.14795274100973, 0.249946445208908, 
    0.356689315482617, 0.259627706023729, 0.190022187971905, 
    0.176066287383826, 0.166150332291291, 0.165461592864083, 
    0.146079170688076, 0.140969512600415, 0.188080726295362, 
    0.190569756537173, 0.128254090326782, 0.142782274976803, 
    0.226189964615704, 0.176677492411692, 0.0971423704208837, 
    0.117040841330136, 0.152645935253262, 0.307174611748126, 
    0.236098819944365, -0.00823983725059692, 0.0814259723307074, 
    0.647820820704013, 0.280158786945738, 0.282593577686498, 
    0.173545707249754, -0.386652164435492, 1.09114053322535, 
    0.712744648820948, 0.580472901576369, 0.872980200175874, 
    0.015942929013061, -0.36664835794605, -0.007525364101083, 
    -0.155757950861245, -0.118168186464786, -0.0680452675818894, 
    -0.24498797570217, -0.0463910715480277, -0.155844869626061, 
    -0.0658198943802684, -0.115231166964164, -0.0684449602011923, 
    0.0248660190444151, -0.211550963575064, -0.0447737653946982, 
    -0.0534078608970565, -0.208364531753816, 0.0684147279830899, 
    0.0421092545834209, 0.14717224288818, -0.0973343443383406, 
    0.140055061865857, 0.0680003012741967, 0.00684445803524329, 
    0.00650948372444947, 0.176657736828844, 0.260247356585653, 
    0.231007141440508, 0.0550627854618887, -0.121682220572665, 
    -0.167951984269208, 0.574707863924844, 0.0972618496262844, 
    -0.270666026121824, 0.0329395665848094, 0.58341839752955, 
    0.197507344484989, 0.103369014131576, -0.137393319012745, 
    0.284629164877512, 0.260376530430373, 0.0794719423652945, 
    0.640549135202382, 0.542094495078762, 0.144866670831394, 
    0.0144603998656582, -0.17722340759401, 0.40330318957957, 
    0.67565272241682, 0.400833666666482, 0.180365560195979, 
    -0.258760310565787, 0.372552074140031, 0.322869373753393, 
    0.132259407624425, 0.53156014621746, 0.343437912814212, 
    0.0529850710418115, 0.404244270933999, 0.445415305513624, 
    0.0314392416064754, -0.263168867913601, 0.111856831915366, 
    0.443329722536664, 0.0221953902530776, -0.107806982794754, 
    0.0887292520994181, 0.181024643217588, 0.0883762206916278, 
    0.203284554159074, -0.0296743494205907, -0.304606681629528, 
    -0.00815361222396115, -0.112055047588388, -0.179071474797415, 
    0.135327422324666, -0.197533582469221, 0.0120551033415937, 
    -0.096316726836317, 0.0106936848725091, -0.22393506353073, 
    -0.015121288759356, 0.0802280251777151, 0.148079117351762, 
    0.172964138406228, 0.164125213612479, 0.174848934856468, 
    0.249315633296385, 0.288364165190277, 0.23271341488144, 
    0.219875743192138, 0.337810191839746, 0.29517734685509, 
    0.201069622690739, 0.367380380592444, 0.474703758156315, 
    0.24692917121176, 0.153595297722356, 0.582642392898723, 
    0.423894376397142, 0.100213197301038,
  0.180615424580681, 0.0610478053803121, -0.0107802864368424, 
    0.109865533685772, 0.108998274879038, 0.0263123181290698, 
    0.0593077771412051, 0.168951829773761, 0.154647095589361, 
    0.0492013804838727, -0.048834290287034, -0.1035464200372, 
    0.052399150431013, -0.0253917769157411, 0.0656601586056578, 
    -0.112082915023077, 0.0618627861270828, -0.193499272218856, 
    -0.0339959530382964, -0.0950105550984585, -0.0603110868406047, 
    0.030376800554068, 0.121198572312205, 0.108763577257946, 
    0.0839179383645975, -0.0456046681843872, 0.142277098626027, 
    0.287269876205467, 0.0352695745694803, -0.0897222257816946, 
    -0.0955838167421926, -0.410050999953509, -0.131642490031024, 
    0.759351378258627, 0.294396994246675, -0.13887413863381, 
    0.171997608384581, 0.556765032030748, 0.247775346949117, 
    0.244409443642486, 0.797863955919515, 0.0815294965344284, 
    -0.00175973551005543, -0.127284513142502, 0.145691152895745, 
    0.305994135258535, 0.337135297657945, 0.268288957545188, 
    0.382416537458286, 0.225069754633463, -0.307846631129495, 
    -0.128981672721171, -0.229178289110316, -0.0328283316100745, 
    -0.265539611142742, -0.143639813784672, -0.00583835504651402, 
    -0.167449940103546, 0.225029518351159, -0.15584605043147, 
    0.155322788922536, -0.0136372994558714, 0.0458371263920635, 
    -0.175370463474783, -0.0333443391781176, 0.00726042733403237, 
    -0.0885617393212099, 0.101889094712047, -0.0432001556366908, 
    0.0542058318014524, -0.0786430645983158, -0.00524226593877422, 
    -0.00131216136964414, 0.02232659517842, -0.104329907415492, 
    0.0244407380813206, -0.0412493168628981, -0.0440049707520533, 
    0.0784146591416185, -0.096867189772247, 0.0167329723787877, 
    -0.00881176303584411, 0.00849839513048123, 0.0212104804535816, 
    0.0155504208681757, -0.0299463577426594, 0.00687348741718782, 
    0.0591406310021825, -0.00881089964111424, 0.153565884720087, 
    0.265395279128324, -0.23674510270084, 0.214405218023687, 
    0.772643450980665, 0.340664378140015, 0.453744658136816, 
    -0.387021955848109, 0.410516359326964, 0.611305669300554, 
    0.0882862853496293, -0.252506639910911, -0.160455328651132, 
    0.464705891908841, 0.333249516916119, 0.119267286800963, 
    -0.179411701882293, -0.0535871478899668, 0.241399814746004, 
    0.565855743284981, 0.110759708176004, -0.284513294809487, 
    -0.168583920175543, -0.225205986340559, -0.112140309790482, 
    -0.225184659891606, -0.148780897999762, -0.0567511309282554, 
    -0.153275719740845, 0.0826292664642486, -0.283815890629661, 
    -0.00530305856975171, 0.19262122547538, 0.0685962119730685, 
    0.1667131436145, 0.362761104460932, 0.210825145877412, 
    0.0287412886336034, 0.350957117888647, 0.474428116022711, 
    0.178034475572591, 0.0304991623191388, 0.0174684245028444, 
    0.0805990600216738, 0.0876621148293727, 0.117416048282623, 
    0.0931163990005052, 0.112892980938518, 0.100348819890827, 
    0.109784015950591, 0.047548189260046, 0.0691693429224909, 
    0.0803181516507014, 0.0989734368299741, 0.168052785447945, 
    0.188931194220909, 0.134809359296699, 0.123312221591804, 
    0.219036300409279, 0.169559400277878, 0.0436177952127668, 
    -0.0336142279252542, 0.316867738747468, 0.420776622752763, 
    0.184059422187447, -0.0763185199723975, 0.485865054374795, 
    0.35137840462271, 0.106179363511562, -0.157037470273928, 
    0.235984349286934, 0.432857693346921, 0.420818767645617, 
    0.164809438565282, -0.209345121602792, 0.0161405064930212, 
    0.677213922154032, -0.0755721409517595, 0.640612374683147, 
    0.784107715162072, -0.15319569100732, -0.136150806445915, 
    -0.085234054502835, -0.0725941640012147, -0.0516901595466795, 
    -0.0558478947570501, -0.0509651358976637, -0.0209115597082542, 
    -0.0710423042760772, -0.182719082908797, -0.0431173344770656, 
    -0.109893307645457, -0.034142826042929, -0.0624434948701695, 
    -0.0891882380528141, -0.00964341138507699, -0.0637496774557937, 
    -0.0833050355645825, 0.0223503775376936, -0.0539758756169842, 
    -0.0312605574271166, 0.0707195675667613, -0.0280714737638799, 
    -0.033803838331921, 0.427337613381076, 0.0868221998807854, 
    -0.0728048011121564, 0.0548418275396206, 0.346123272448628, 
    0.0670275544820212, 0.174379296087751, 0.503625676448803, 
    -0.360470683860489, 0.379739894292712, 0.899425588780207, 
    0.656822390973594, 0.234192463623177, 0.0340756679435958, 
    -0.518055063992497, 1.1202760679072, 0.547900201131993, 
    0.312879504199861, 0.265913552208245, -0.159357735175104, 
    -0.147666509077894, 0.129007313828438, 0.262187071687487, 
    0.583926783236883, 0.358425103669116, -0.0199617576209801, 
    0.375347723469098, 0.407066051197069, 0.0856127262428266, 
    0.084211303153586, 0.22848759098192, -0.19414400647949, 
    0.240509878248239, 0.441407325186476, -0.0882670502443569, 
    -0.0668157336531006, 0.130826118809099, -0.147347495155256, 
    0.190159773427329, 0.188237989464487, 0.299511782748352, 
    0.620530426423085, 0.251329351637224, 0.12575593789773, 
    0.405175850315902, 0.0675855064410397, -0.0583178654062787, 
    -0.012530746271412, -0.139641379594134, -0.0159340328309868, 
    -0.141903603712448, -0.0613055877163778, -0.0995601268300888, 
    -0.0906129118006534, -0.0782910491988053, -0.00951832656681023, 
    -0.145324319926833, 0.0489023144701035, 0.0640610475003977, 
    0.0795254072634785, 0.209600007970868, 0.138991503808382, 
    0.0435387438104497, 0.299264170374131, 0.13957830060905, 
    -0.0450015225618665, 0.113019766177555, 0.700327990585298, 
    -0.187853014628336, -0.0883058242968236, -0.100906092677265, 
    0.702438311535576, 0.0214174169596151, -0.154641687885727, 
    0.263403504406143, -0.34082502365531, 0.939063102223145, 
    0.677833952083656, -0.165001899671179, -0.0405083610570745, 
    -0.458126649963994, 0.0445050428725926, 0.25330877716215, 
    -0.065584654612686, 0.260731557475675, 0.227215623829294, 
    -0.128239019894022, -0.0450333662689953, -0.241532916299389, 
    -0.00487580036740154, -0.279079358319142, -0.0878134898563528, 
    -0.152890635736417, -0.0713105335223419, -0.0371894502011475, 
    0.219303739009393, -0.266588186432587, 0.0323520147025861, 
    0.303111673244237, 0.146980077005324, 0.0649173525457919, 
    0.120696775158462, -0.087534969057084, 0.0917613050977515, 
    0.738957225731601, 0.179465779081936, 0.227740568317053, 
    -0.515846502077048, 0.324179640574747, 0.660037097850268, 
    0.0924554560623978, 0.0598720770975893, -0.334550036914175, 
    0.672034113897303, 0.432926009139982, 0.210451539898071, 
    -0.0325069064737598, 0.339609104595543, 0.428764029215998, 
    0.197705098699903, -0.0523625146784134, 0.234248940597351, 
    0.289997146330648, 0.334053272996778, 0.231224446243181, 
    -0.148133065928865, 0.026292653492955, 0.642325835882623, 
    0.173994302602168, 0.102284177909632, -0.0179984560037926, 
    0.494161153242338, -0.0409527857878347, -0.217840030153532, 
    0.0397654119448743, 0.407767380940024, -0.0142167403036819, 
    -0.119635584414488, 0.16406788739409, 0.265175388892688, 
    0.0242951599159578, 0.0834713471525109, 0.069772085948426, 
    0.249804584840612, -0.0794165367290186, 0.279193722266691, 
    0.408021986612423, 0.047227975424496, 0.0164191676742873, 
    -0.0198957765109733, 0.134195905019841, 0.175508231036757, 
    0.0902336765956197, -0.00161498126739204, 0.237242305397684, 
    0.12903384308345, -0.0876940348778044, -0.0862996768092198, 
    0.156100443956207, 0.475525602869428, 0.283643887213328, 
    0.107243812606112, 0.498756626229819, 0.28863183144311, 
    0.0831028353008557, 0.0469301528726059, 0.445138035751203,
  -0.0323481050834985, -0.0852079388530309, -0.0724474099771218, 
    -0.131966440923083, 0.128474420694986, -0.00778375659664693, 
    0.0583519128023379, 0.123684937354556, -0.0852330312451837, 
    -0.0644913313901314, 0.0016515674766838, 0.0162452153176108, 
    0.00568389509237446, 0.0168119607580009, 0.00749741000847372, 
    0.0242785655893198, 0.00620106720311847, 0.00300185031979947, 
    0.0804481399130724, 0.146140133064205, -0.0417900807303719, 
    0.0856468094056788, 0.339788373870631, 0.396981299803382, 
    0.261930929981987, 0.0254047225032624, -0.0597947636134404, 
    -0.310858344699835, 0.581554366429034, 0.303778524595724, 
    0.0716580086025282, 0.331700761385456, 0.23653972573655, 
    0.116961270891655, 0.151787184855812, 0.0267996051812708, 
    0.123974062069114, 0.503283499050565, 0.181231031935999, 
    0.00826423460535669, -0.0459358706150708, -0.254750882880582, 
    0.0604834901094055, -0.101535801517955, 0.0528991421516625, 
    -0.153129946839013, 0.041356721312638, -0.182849220302032, 
    -0.0463107100404443, -0.20186050551837, -0.148605974994076, 
    0.105356637278683, 0.157948867035046, 0.0347190871024092, 
    -0.0659574078367003, 0.292101388313562, 0.226031238415944, 
    0.043491764994728, 0.133794159974807, -0.355134242137124, 
    0.529596263402357, 0.308073761116946, 0.0882317735315034, 
    0.0841878115547058, -0.374550913446359, 0.21994231453744, 
    0.615768031145945, 0.420958504143165, 0.251548827862866, 
    0.0912576971540014, -0.190478836474092, 0.0196427273733811, 
    0.210562961722218, 0.478189241660193, 0.152571502269491, 
    -0.115955664736396, 0.185605799297895, 0.0797292581636777, 
    -0.21303602642882, -0.039679489700485, -0.323758054862312, 
    -0.126023807836907, -0.243039945514792, -0.087379740808283, 
    -0.291105363987199, -0.106228317620244, -0.185087195764854, 
    -0.212861056467668, -0.0102029593582775, -0.201696525956905, 
    -0.0180921616723179, 0.0550766814294082, 0.0122981468722212, 
    0.0325947625688692, 0.0414998151795352, 0.0445851026690486, 
    -0.019250755394253, 0.040899011699683, -0.0183900753401305, 
    -0.0341067514588629, 0.0390821434078331, 0.109803698009639, 
    0.128675712165115, 0.134553955792032, 0.142111988512277, 
    0.0802106936335443, 0.157260589586997, 0.402013793054013, 
    0.0583428273560068, -0.176251957096237, -0.152931001812226, 
    0.198191680323909, 0.61474304066597, 0.35182806571013, 
    -0.0903616030157814, 0.528668673260825, 0.484842951160587, 
    0.163543148793169, 0.111742806685875, 0.510478445487006, 
    0.156415125223095, -0.00672777109290204, 0.340914931485206, 
    0.323219753775777, 0.0674701544456689, -0.303618655377682, 
    0.113898240146194, 0.37988667821229, 0.353628802868149, 
    0.101872151604016, -0.178270720003947, 0.0584027773123573, 
    -0.19196035442076, -0.0436122817058929, -0.409784063570022, 
    -0.0842035433669629, -0.132579189724201, 0.0609972116012795, 
    0.222232593118203, -0.431276256570349, -0.163813336008534, 
    0.219456643901604, 0.0534073039195161, -0.100300962774444, 
    -0.0404132791171394, 0.213132026918867, 0.231600580425711, 
    0.370379331405073, 0.434222588293323, 0.0309084473468217, 
    -0.321700661067154, -0.0537228878037913, 0.857353260538933, 
    -0.123540171283885, -0.0764433858917738, -0.421610537411823, 
    0.810679241146451, 0.395901163123085, 0.085129988217715, 
    0.79599046763008, 0.401136574850838, 0.038741622909876, 
    0.225176531191047, 0.735401946567437, -0.163089480468522, 
    -0.275545761028437, 0.113230282132156, 0.404302369750039, 
    0.0755822349606428, 0.31740649164951, 0.37450467359338, 
    -0.0974100410827974, -0.113217758145367, 0.0135784132139865, 
    0.240512409581837, -0.0212139669249001, -0.239422210679448, 
    0.00643715413551359, 0.258932719208003, 0.057095642565321, 
    0.00681135414941477, -0.046183583275592, 0.141716606253278, 
    0.246059072118367, 0.140128927541557, 0.0513449698346071, 
    0.0752696769361099, 0.243180338177701, 0.0680109461006602, 
    -0.187558730259886, 0.0289173067247357, 0.451352175010799, 
    0.117847931473501, 0.0795812608111282, -0.210483580720886, 
    0.446888556850154, 0.272156822367753, -0.0519204829935346, 
    0.200831248531345, 0.530888769480536, 0.162811169183026, 
    0.127159966740331, -0.0286068469870303, 0.260076078822033, 
    0.179578330896961, 0.0814545727421862, -0.0234946140646831, 
    0.491822205486776, 0.0234271443383673, -0.113808146785784, 
    -0.0611151094120213, -0.231384671377075, 0.086724695124282, 
    -0.139843731755728, 0.0833482313914309, -0.231397031694804, 
    0.0600210645735884, -0.165039167875556, 0.0310977029311251, 
    -0.270797318608895, -0.0396616908071154, 0.0524043050445047, 
    0.16287311085457, 0.197156811699102, 0.150161077125363, 
    0.100252847566407, 0.182924283170723, 0.309667009415815, 
    0.274366673917997, 0.256633204094572, 0.308455467379629, 
    0.169891986354042, 0.066175100982119, 0.554723365241324, 
    0.543423129510152, 0.182023047486406, -0.0764447962752714, 
    0.525069262523747, 0.53587944049019, 0.161378996482694, 
    0.0456138170332196, -0.216033891714644, 0.226672233263771, 
    0.548465480928887, 0.330721005537763, 0.113923724715559, 
    -0.0258332623371419, -0.00629088824883366, 0.745425098419965, 
    -0.000600617708291056, -0.0581882714830609, 0.0179111321589245, 
    -0.0951966602176225, 0.649681531082331, -0.0541183750175449, 
    0.0578366994374624, 0.431359652283093, -0.0197697576738947, 
    0.509183930349269, 0.0145535998384209, -0.248432910213712, 
    -0.0339146745478509, -0.448658217828256, -0.136378757102646, 
    0.0386433956670427, -0.36774912740609, 0.121469882870628, 
    -0.115242310172629, -0.0305123211092589, -0.345800884709748, 
    -0.104981619489539, 0.0818080863714222, 0.140654558287294, 
    0.221210383687165, 0.188679188490813, 0.0869563448670498, 
    0.0515796892644561, 0.190287929420994, 0.220387948316296, 
    0.154233307741183, 0.144347677521513, 0.152419600143718, 
    0.164036456248271, 0.193164066396107, 0.209481239398843, 
    0.15594099037303, 0.139318767614623, 0.290646495800816, 
    0.221844639485363, 0.125133865628776, 0.278551042755416, 0.1692075677688, 
    -0.190766748496948, 0.579110593062302, 0.417647061438321, 
    0.0115909956971189, 0.00920436416913354, -0.302958469545396, 
    0.153185339475132, 0.492156526373429, 0.126798046636462, 
    -0.0192595710406216, 0.413050471809276, 0.0683109051217015, 
    -0.121498080713192, 0.11089990158212, -0.292454631448174, 
    0.0969336213924978, 0.234017238510388, -0.0242043594976972, 
    -0.0778583282793577, -0.213742959410401, 0.0818176363374163, 
    -0.0709719699093815, 0.082744547353484, -0.17517145366188, 
    0.0811869584618188, -0.0761001995328982, 0.065437640890942, 
    -0.297234527745495, -0.0545308932527478, 0.115808441049201, 
    0.142063756491032, 0.088650270908793, 0.0877124015654449, 
    0.124464241409852, 0.238690417585259, 0.383105276995671, 
    0.285062571059235, 0.104419364919425, -0.167605338364795, 
    0.323439167877746, 0.673404296485302, 0.176608366660728, 
    -0.301148319297353, 0.281678800677662, 0.742026745140103, 
    0.0544445593145392, -0.272183186273762, 0.075723964355153, 
    0.631250484882148, 0.150284930406036, 0.0217215180380139, 
    -0.169321407281947, -0.0471241338492771, 0.7270615646865, 
    0.211671029034541, -0.160578166220784, 0.172898374570079, 
    0.597119684702349, 0.0489722011897862, -0.364235276151346, 
    0.241231580266525, 0.364811612680183, -0.0404332028878641, 
    0.0333162794218874, 0.19249540075442, -0.132008968471335, 
    -0.12428312363898, 0.542052602814199,
  0.555816613731774, 0.236888192472709, 0.0138307042804144, 
    0.524365260978282, 0.314155265086601, -0.0599560985841355, 
    0.752342153962837, 0.617978301504055, 0.187076205081639, 
    0.178488555545018, 0.591572268879677, 0.372327781945025, 
    -0.0422587272891534, -0.339600455126574, -0.417427492725962, 
    0.493958934323065, 0.402915134646624, 0.18568044395328, 
    0.164769999497388, 0.204153098843472, -0.189334088919801, 
    -0.359469205665467, -0.113941441412227, -0.270646760948633, 
    -0.0828730268792755, -0.285912247782318, -0.153421865435186, 
    -0.137492579914489, -0.253730619931641, -0.0374320645147903, 
    -0.112156319338071, 0.137905300054864, -0.109850152580975, 
    0.0578671220787226, -0.170372815248526, -0.047686504687146, 
    -0.025263241418117, -0.0991203925111115, 0.0521440700292709, 
    -0.0971278876892256, -0.00988001708835203, 0.0677023643947446, 
    0.105102913338313, 0.114977280131967, 0.123540881790707, 
    0.128933299575238, 0.130241066827834, 0.126514224843237, 
    0.113634626685546, 0.116328183799919, 0.15830405423562, 
    0.157043735874624, 0.15230879262562, 0.169610476709295, 
    0.178320301012246, 0.145724773696565, 0.133506554179802, 
    0.196234747994718, 0.196729320448022, 0.106130448327727, 
    0.065808395623861, 0.252939631068006, 0.285408122445414, 
    0.125070658901735, 0.109525271933498, 0.356287082592262, 
    0.269681256384107, 0.151034723173144, 0.116832755256024, 
    0.113070974989844, 0.695284420841333, 0.343567692571172, 
    -0.111636223753961, 0.206358082570626, 0.626509393111135, 
    0.27067902328947, 0.12078117442601, 0.19510688936586, 
    0.00203592079982084, 0.62481128469131, 0.327549261929099, 
    -0.0631510920255997, -0.0776968118634789, 0.0290697314803671, 
    -0.0893274862825962, 0.035819463058947, -0.0011081166463336, 
    0.150559888425702, -0.0174179095882009, -0.158752959819811, 
    -0.225484667604056, 0.0446204763778278, -0.180017771599022, 
    -0.0333350684931403, -0.117845008123722, -0.0255766838247589, 
    -0.216374115324606, -0.0916528673391719, 0.0607468114232411, 
    -0.297956174941341, 0.112199197526889, 0.115558986453904, 
    -0.0650883597462578, 0.0771079031287903, 0.212206522704289, 
    0.355069743267134, 0.232044484919935, -0.0500972473152992, 
    0.354817965261855, 0.0661628434270645, -0.0310943810630439, 
    -0.0330189757615051, -0.41139291672557, 0.877303796960914, 
    0.35369981705512, -0.137273786619999, 0.147953468999829, 
    0.72132079512915, 0.354925466414816, 0.104537737825388, 
    0.177714961419356, 0.421324064110919, 0.308890039809562, 
    0.0834524014358458, 0.308010386473673, 0.533458327223381, 
    -0.0196133690207174, -0.157216326443765, 0.14917094661555, 
    0.312811747559774, -0.0674991992999101, -0.00643770075416659, 
    -0.0899736661983319, 0.0647753048691766, -0.0873529228326413, 
    0.151081422685346, 0.00375173951025758, -0.0261399890592064, 
    -0.0601070548482133, -0.0965916555268703, -0.196469548360835, 
    0.115651029579982, -0.178150403148905, 0.0183990252105941, 
    -0.167926756598192, -0.0133425170529197, -0.173812270341028, 
    -0.0829490618812373, -0.0176472986402904, -0.125894801445256, 
    0.0812663104229365, -0.0707465493525999, 0.0317744385857506, 
    -0.0516413943844593, 0.0291467530519803, -0.087323601562382, 
    0.0175342402177089, -0.0476747867097761, 0.0223839261384845, 
    -0.0947749641604353, 0.0175954016653996, 0.0497286698097043, 
    0.0637282217135915, 0.102576821404901, 0.11839958546588, 
    0.0795827502641332, 0.0895368901950251, 0.185223856885135, 
    0.0885097042173019, -0.0344763205883697, 0.0634776590312031, 
    0.161735055135955, 0.0924198011857074, 0.645922500137748, 
    0.347525881541208, -0.00470079725095839, -0.332503008463695, 
    0.0711547205557154, 0.587802766284315, 0.52415880364357, 
    0.156295624220079, -0.263086816689251, 0.0912474212840984, 
    0.413093870582774, 0.213831077921099, 0.316593448227957, 
    0.43058843005632, 0.318598063329544, 0.771794579381969, 
    0.0529659675438442, -0.286504429980692, -0.1101794631467, 
    -0.115745146910183, -0.0811254476268017, -0.173963226635468, 
    -0.0997729720394371, -0.185848249096573, -0.0973575320823043, 
    -0.136481791922257, -0.183428740262156, 0.0288893985074962, 
    0.0185647532128926, 0.0657630851427114, -0.00870582134537205, 
    0.0402042414636425, -0.053022769736009, 0.00593197150484516, 
    -0.00382998382073468, 0.00834354355766198, -0.00248370512032126, 
    -0.0779182949698494, 0.220792385563701, 0.249530491671853, 
    0.0660404107557359, 0.157724870326775, 0.278427493747583, 
    0.53424134087692, 0.288494426587039, -0.101391599162998, 
    0.447768375074547, 0.193566344347856, -0.228213762432254, 
    0.018545133920425, -0.178883810367721, 0.415713029371564, 
    0.254535840239534, 0.0291542127944477, 0.188531110058681, 
    0.678243009308656, 0.130835273512539, -0.0568223973119358, 
    -0.176733406337711, 0.110350647892083, -0.0237480265064873, 
    0.0715358735115587, -0.0971935728945766, 0.0905522577365656, 
    -0.0836680461962464, 0.104825791142173, -0.0873142357175893, 
    0.228904732813673, 0.0265935524470673, -0.0921659050069575, 
    0.315630094009298, 0.496519017034431, 0.14016821399651, 
    -0.258950678308775, 0.271549973313698, 0.479158090872781, 
    -0.269987693662255, 0.276979332606311, 0.853895369802279, 
    0.110900509185899, 0.126615706800632, 0.227919506412511, 
    0.950450053331489, -0.086550237018607, -0.0358954478522115, 
    0.0579834102052331, -0.0896754606224773, 0.124367967228635, 
    0.951911537497545, 0.315277521396614, -0.0630631309001125, 
    -0.321931530734941, -0.188666086055572, 0.297132515082433, 
    0.61924380451014, 0.360908015744666, 0.21868534907759, 0.368754622787627, 
    0.00580963127700807, -0.124827955182014, -0.297767750379228, 
    -0.230507019636497, 0.416344264267413, -0.129380917130759, 
    -0.172649743983478, 0.152927869844059, -0.00732131804277202, 
    -0.224723791309764, 0.0713735041297693, -0.231334796554893, 
    -0.0809405331040561, -0.153560991146224, -0.12737805335148, 
    -0.0647466605088655, -0.141141379857299, 0.0577057259766738, 
    -0.104512279005938, 0.253544097641514, -0.0297755259676031, 
    0.0509100207688189, 0.386480911086845, 0.208240909907107, 
    0.0607813601701764, -0.0300868553836957, 0.0417707487721207, 
    0.379781991190063, 0.466797951504841, 0.192910617556393, 
    -0.347947331309812, 0.128076630159146, 0.572631489414756, 
    0.177577351163769, 0.0518353330944718, -0.149416623272592, 
    -0.135479240735878, 0.444308799565706, 0.423876028613666, 
    0.224029206067304, 0.229727644691425, 0.160305962031729, 
    0.00804081006153609, 0.243567763881023, 0.466219000700378, 
    0.265515243072418, 0.101030111015426, 0.00116507171195274, 
    0.140807241479756, 0.293795278841626, 0.364016734861796, 
    0.362559002600064, 0.174282794602767, 0.0174382582593906, 
    -0.00561410206415174, 0.0655399353270327, 0.138682144783005, 
    0.665419082983105, 0.404902804266458, -0.0545948838492706, 
    -0.175969321852353, -0.0302724134483466, 0.59796127385897, 
    -0.053933027744463, 0.0493523446396161, -0.084031506090015, 
    0.238406814207093, 0.264526218439645, -0.134998058187779, 
    -0.17638367950194, 0.00763559175417901, -0.350642374459603, 
    -0.079693147068383, -0.156218757132654, -0.246229795165718, 
    -0.00497263299122559, -0.115028667707845, -0.0050485551433984, 
    -0.222252566706831, -0.0328922531219192, 0.0926947608708035, 
    0.0885920607586834, 0.0976553263336393, 0.20088643846895, 
    0.241895051070506, 0.226597203338132, 0.142005296724022, 
    -0.0575774611178805, 0.164141150930396,
  -0.0991349422147062, -0.136856569183568, 0.0179077644946602, 
    0.00460227325353964, -0.0289842720576024, -0.0254985639271302, 
    0.0410719036961252, -0.0862338949033952, -0.0358698560357523, 
    -0.0991530450252194, 0.0860512244541838, 0.0689728593466628, 
    0.0498765296958439, 0.0426084107756637, 0.0314254140199264, 
    0.0504863754040509, 0.114736410050232, 0.0486111445152888, 
    0.0484863826237199, 0.0491119671485885, 0.00820111917406718, 
    -0.0248128551525644, 0.0121207293721973, 0.0345114619927824, 
    0.05108662092573, 0.0131149408043378, 0.0590145534690197, 
    0.0297785610034366, 0.0663018012441974, -0.0548988007054229, 
    0.0335708215095601, 0.181006485312004, 0.134035891938903, 
    0.00981950260036069, 0.0748081631578684, 0.290914518605113, 
    0.298241170701558, 0.11902608266653, -0.215609808775619, 
    0.169635571337153, 0.463084404047621, -0.0786790768460184, 
    0.238612566216301, 0.716971246018329, 0.115898615520625, 
    0.0402566834034577, -0.00467816778585738, 0.743449042682191, 
    -0.0244203553653992, -0.204299615902484, 0.161353755319419, 
    0.26585653887855, -0.0883377164074409, 0.00916408734361859, 
    -0.0669594742332436, 0.154838855512837, 0.0797210672499237, 
    0.287504698058343, 0.12638672076356, -0.17235468352096, 
    -0.221817683127195, -0.025533751871544, -0.291031636392469, 
    -0.175409454019727, 0.0698794010691798, -0.163057499231996, 
    0.0709721450821638, -0.0231629054607691, 0.0965808086355039, 
    -0.249336469631434, 0.0814456013179338, 0.101586921229049, 
    -0.00987720388334774, 0.162562325771557, 0.312157386684436, 
    0.165892658581302, 0.0404839342835785, 0.105731258753902, 
    0.300303072227551, 0.378786457461663, 0.235490435101788, 
    -0.145804211492777, 0.122614178656406, 0.761837064887407, 
    0.280946633904293, 0.0484933672346428, 0.0646055118690811, 
    -0.130721593304263, 0.648339109127768, 0.708238430440064, 
    0.157542363403587, -0.044733832686219, -0.332109787388819, 
    -0.265461642342002, 0.567409530456205, 0.164510126047656, 
    0.145498929684477, 0.314706733047733, -0.376225799113747, 
    -0.200696513661603, -0.275711395810503, 0.0312770677614223, 
    -0.248206005210967, -0.033042355188142, -0.313790848700717, 
    -0.158582812879392, -0.0785385047126373, -0.247473073646813, 
    0.0863551405757826, -0.198516101331751, 0.14981893280199, 
    -0.0299143666312508, 0.0836093400109189, -0.000648651600946987, 
    0.0758769405090677, -0.0226909819579066, 0.0699204626935412, 
    0.00682367350196751, 0.0408767454499614, -0.133259196680386, 
    -0.0261287697046485, -0.0365249797800447, -0.0438231397207704, 
    -0.0350904053587674, -0.0236807353113463, -0.0331401490662035, 
    -0.0416377554476531, 0.0770989429664215, -0.0614847146689138, 
    -0.209147731098222, -0.26035383222524, 0.169300181712081, 
    0.406850817875136, 0.166327614802264, 0.248019510589272, 
    0.0746289249281851, 0.615466101387645, 1.10940735042043, 
    0.117494480330367, -0.122617166359894, -0.244837201944885, 
    0.400964720378249, 0.439056458744698, 0.283404073432134, 
    0.18052567937853, -0.391818393604193, 0.48858823404316, 
    0.671351514240644, 0.224065992601777, 0.0777862495209393, 
    0.275994130084094, 0.267983693163229, 0.0933811765553314, 
    0.0387484921023714, 0.0197623226366471, -0.00140413184295488, 
    0.0187219814081333, 0.0697047532858931, 0.0473697322404653, 
    0.0508357893991427, 0.0101341401891356, 0.135179687009228, 
    0.157303927095635, -0.178975152522443, 0.335654544287383, 
    0.636454796712306, 0.24338411151387, 0.0235761256477917, 
    0.58048650101016, 0.240585180446042, -0.00527523948278816, 
    -0.0166330881185306, 0.0758895858702995, 0.0642357785520577, 
    0.133973838937587, 0.155833556752608, 0.0630487653089228, 
    0.0330843017771393, 0.0269296259041621, 0.0269940190459998, 
    0.0116639806581039, -0.0966907451155682, 0.0652587217242838, 
    -0.144014163713216, -0.0161452684281061, -0.153334808430586, 
    -0.049127108757858, -0.0581404049209936, 0.0817903463860452, 
    -0.130262426051643, 0.083682300478744, 0.09610434359771, 
    0.0523244545581494, 0.0986567030474613, -0.00458597020583618, 
    0.165613188986264, 0.24072649940581, 0.0449655425799662, 
    0.114195662646303, 0.220006946697483, 0.136258608412045, 
    -0.47205692737175, 0.507302501877231, 0.540891670670739, 
    0.356103742694018, 0.584438590253401, 0.252298111815092, 
    0.24987834162122, 1.25852340908321, 0.181203853340532, 
    -0.144014051803833, -0.198362113584099, 0.0428344167331837, 
    0.172342284800198, -0.0988750292788953, -0.125338888467834, 
    -0.0356290770849452, 0.224141536647621, -0.0360834400539648, 
    -0.0354434387434925, -0.186380257348644, -0.192093917045713, 
    -0.0728129434136911, -0.243953941420345, -0.155737977867237, 
    -0.169290553714357, -0.178087206915255, -0.100441997424552, 
    -0.0758856465549858, -0.163577209481807, 0.112686074274574, 
    -0.0818561755142167, 0.0754816188996938, -0.0693147843469975, 
    0.0511789416154093, -0.119381856202212, 0.0377572808958122, 
    -0.0586722313001487, 0.0446855404813427, -0.177603440429977, 
    -0.00829917006874173, 0.0634902768999748, 0.06223112468171, 
    0.074416554225583, 0.126325668904296, 0.124809399788754, 
    0.131222519273258, 0.186411883857009, 0.119918520570035, 
    -0.0436965450710287, 0.173587278784568, 0.390042628092734, 
    0.173253063209111, -0.0841508918318218, 0.171216836089641, 
    0.521414710749703, 0.348725369154771, 0.169364069716835, 
    -0.209598685712508, 0.432254559710321, 0.427408205245031, 
    0.0992121794920026, 0.00813049264672446, 0.553661622046391, 
    0.386032224549766, 0.0817246915472554, -0.295931670924417, 
    -0.115678730470285, 0.505073748630424, 0.302731171574178, 
    0.268368365464005, 0.319517654465346, -0.15309017015615, 
    -0.287242388484639, -0.00445949681103136, 0.175976366238256, 
    0.13957145401215, 0.294462246228834, -0.034376362143313, 
    -0.180954102574147, -0.208888497018263, -0.0502117062795629, 
    -0.255406746172463, -0.160260850675371, 0.0918899422044032, 
    -0.220086263437291, 0.111586574209412, -0.0770445783517498, 
    0.0684429959058388, -0.256749300268839, 0.0353471435663993, 
    0.0804329134360319, 0.0197043015876541, 0.152647861070366, 
    0.283283537544512, 0.16799312376822, 0.0745536392164748, 
    0.244285056187906, 0.267842077397566, 0.0975877277201788, 
    0.0838681465108818, 0.392294392940671, 0.591204152690101, 
    0.342218280339073, 0.0996749044032569, -0.211602947829863, 
    0.722905564203349, 0.693429897328596, 0.205176977839468, 
    -0.370261389081404, 0.468698885927843, 0.510850409587746, 
    0.207225609692885, 0.184173629763101, -0.175825686172742, 
    0.590180612801304, 0.16010847339292, -0.101077060594796, 
    0.0691484568953346, 0.669493896727338, 0.0249627408835018, 
    0.0185207296444023, 0.0130167458832745, -0.0370141800899695, 
    -0.00095547236288171, 0.140734529965201, 0.0385034842218203, 
    0.301626561042485, 0.114289825850919, -0.0680588062938308, 
    -0.0275122142783661, -0.0802136300209177, 0.00100696433719276, 
    -0.102686018206272, -0.0540167623421959, -0.0250449073521608, 
    -0.0943860584126345, -0.0130561524758115, 0.0564758038594363, 
    -0.101865704212024, 0.193638055869811, 0.0883587400232983, 
    0.481909823906982, 0.265911718648473, 0.0742872831530581, 
    0.0203719821202754, -0.0429685478069397, 0.634765864883026, 
    0.125980368786462, -0.0498484480946919, -0.320138206006725, 
    0.817613558530904, 0.300884423470725, -0.219490567282235, 
    0.636659747886436, 0.509455000899951, -0.232026836501611, 
    -0.0457355375326214, 1.05773601058047, -0.0326834596067817,
  -0.0313062458409988, 0.0602577319408572, 0.0837077404416683, 
    0.185700485871945, 0.185153202406049, 0.114993192601519, 
    0.146136696460173, 0.15261449924272, 0.0148438996459896, 
    0.272838798794701, 0.359699550760378, 0.0422303907747771, 
    0.27735781550489, 0.453834421213764, 0.136648849904236, 
    0.100419083886956, 0.60015087124856, 0.344446947455196, 
    0.128903591167594, 0.0301789829714832, -0.0209019088688803, 
    0.210181157111444, 0.334084454654854, 0.294305256210552, 
    0.237370760844203, 0.194900853666183, 0.178957181725531, 
    0.193914297583739, 0.207460616846982, 0.221826670038664, 
    0.215922788556101, 0.147265909140569, 0.110520628864883, 
    0.290735130864462, 0.253441279653085, 0.0573355602564412, 
    0.119029888934478, 0.406201561548921, 0.198889129352308, 
    0.157895550474283, -0.151213211522177, 0.405932743857706, 
    0.318853797914534, 0.135300568122441, 0.0786703873414053, 
    -0.136526455775286, -0.0361912380053155, 0.74925398579943, 
    0.241837453164064, -0.0200593789757586, 0.131763528960543, 
    0.309506522463909, 0.125437994792984, 0.359701178674591, 
    0.408093432731202, 0.0851422393996275, -0.0527245723562612, 
    0.53859315311993, 0.161487583098525, 0.000984494859530865, 
    -0.191846228377038, 0.0208926837530529, -0.134451529870466, 
    -0.00628857852450381, -0.0899294911443649, 0.00535691758041394, 
    -0.215029567191987, -0.0659825660407035, -0.0610578966022969, 
    -0.182278558373879, -0.0017642410438416, 0.184082215982225, 
    0.0864654085035021, -0.0157355892446117, 0.366742828065147, 
    0.238201542129335, 0.060093163965769, 0.0429590376734172, 
    -0.220523753642044, 0.187278687247939, 0.40718147324651, 
    0.375570551915627, 0.307081653999836, -0.13068263278255, 
    0.600913288264025, 0.525228865434675, 0.188209957206073, 
    -0.28555112869826, 0.277373606495897, 0.522441857062683, 
    0.0186867787626704, -0.0974349704260516, 0.236124194049142, 
    0.0500025811093394, 0.0140040828984528, -0.0645760023168484, 
    0.110558587929141, -0.152974100389389, -0.361251462676846, 
    -0.112567190874602, -0.222676119047159, -0.232932316040429, 
    0.106410584323591, -0.188146313779494, 0.200601401312361, 
    -0.189754576053819, 0.0920342490433618, -0.0631667756848261, 
    0.105962071971754, -0.26120389076426, 0.00643416010529311, 
    0.0692806616263161, 0.0943592566125465, 0.074678948030018, 
    0.0834548178434902, 0.0507785350164092, 0.0595294851231444, 
    0.0913391341426457, 0.0945327476902958, 0.0379405187684873, 
    0.0788880650737461, 0.108765171499193, 0.122768617826132, 
    0.129318806118056, 0.129048437710478, 0.11300840758057, 
    0.125966605186986, 0.189583000900493, 0.144473060255869, 
    0.0538462620619074, -0.0772035397823718, 0.172379895734605, 
    0.37505326123489, 0.214250944619652, 0.0996511308363026, 
    0.0581458247804261, -0.0911340000192651, 0.271119545529969, 
    0.62634015860878, 0.113368584844997, -0.034267715757502, 
    -0.285790398772466, 0.179539422688497, 0.531198684775039, 
    0.516430394102325, 0.328435640183081, -0.171631722212684, 
    0.722113823152497, 0.419009378842382, 0.0870963571792288, 
    -0.15362997426639, 0.13471006123749, -0.222358841121265, 
    0.109562899948336, -0.274629205566371, 0.0180374146103568, 
    -0.271157062099092, -0.08963221384879, -0.150790059858037, 
    -0.196354143064225, 0.0270840815128254, 0.129651547666046, 
    0.0594278398639516, 0.0869342434170746, 0.146684870107091, 
    0.0890179336964395, 0.0984227251077136, 0.150696869009664, 
    0.140675472629162, 0.0886615658458426, 0.0914675143680323, 
    0.114515826356152, 0.126137728469191, 0.145512041487048, 
    0.170850141159109, 0.122034079473329, 0.0762382761168198, 
    0.253934049245326, 0.160984508096083, -0.0386784982572683, 
    0.195530724572407, 0.322131650269289, 0.0610711293812113, 
    0.340630988826726, 0.299863390005069, 0.231679133390642, 
    0.686780792662897, 0.467756315843716, 0.198462451695771, 
    0.151382425312798, -0.0468312934570871, 0.369031571590918, 
    0.364278888887762, 0.669478063323717, 0.286246539484304, 
    -0.224565099563867, -0.0454120483290203, -0.0728703292842541, 
    0.549905678112438, -0.119251170280376, -0.154676405993113, 
    -0.0426839103112526, -0.0823687959526252, -0.110497308603561, 
    0.0397805448468718, -0.107862008009243, 0.0205571383659292, 
    -0.0451595578179526, 0.059914064094211, -0.142811411901844, 
    0.0452832485699846, 0.122976486714132, 0.19756643338164, 
    0.258847192825357, 0.192774785179226, 0.0721839540183541, 
    0.230768359717469, 0.485113725514424, 0.31539020265417, 
    0.154277228443303, 0.378954515078381, 0.391870612946186, 
    0.0712027739514762, 0.226528109623113, 0.802983200669444, 
    0.298003240207507, -0.00543367732679154, -0.0137726550409068, 
    0.64477719751523, 0.325515681066968, 0.0612967033178526, 
    -0.121879676432216, -0.0208486999016652, 0.381573874109807, 
    0.513203621152421, 0.25323835359421, -0.102445933254432, 
    0.466115722352205, 0.295967654811745, 0.039012942936845, 
    0.272627564406838, 0.340444103214479, 0.263059820180083, 
    0.175082511693058, -0.0271316039184927, -0.0296529603146142, 
    0.00432939116493016, 0.659962275508584, -0.00757414650363134, 
    -0.049217886023588, -0.179167686422123, -0.123802947297585, 
    -0.140450668497524, -0.142327759647991, -0.124244225592218, 
    -0.135381179953684, -0.126897480301746, -0.120723159858789, 
    -0.0389993554268615, -0.17091206146276, 0.0745844958271454, 
    0.0158747829995328, 0.0550823835044517, 0.0358124430819891, 
    0.0547519044795367, 0.0178953078827766, 0.0433909838451672, 
    0.0648447981744792, 0.0576890351770103, -0.0198516520522064, 
    -0.00417869482403914, 0.165752380736333, 0.155987708789623, 
    0.0379567128702702, 0.210367611517022, 0.251047377069633, 
    0.0875751541127557, 0.0144522045623897, 0.00740787294197064, 
    -0.145947980495097, 0.528093757199976, 0.345575412744827, 
    0.139893325496645, -0.160803968579005, 0.256040857249706, 
    0.129774059863109, 0.300403836540955, 0.787990015821951, 
    0.334960097296997, 0.0740825250642742, -0.298479772581388, 
    0.172339700046923, -0.132878384940131, 0.034505862568564, 
    -0.120390705703109, 2.58586835974878e-05, -0.471395890369715, 
    -0.086858546141931, -0.0865058406507222, -0.359317881721547, 
    0.172283756516194, -0.0482943680621815, 0.0484971005532222, 
    0.0507160474718551, 0.0348087839880927, -0.0926049052140089, 
    0.0632059000122598, -0.0634045100591736, -0.00309211588070082, 
    -0.105056110309815, -0.0712533953047074, 0.0283891361232057, 
    0.031479386681297, 0.010312826688019, 0.04494653440962, 
    0.0511008593595058, 0.0452305855808919, 0.0799930032969985, 
    0.0685382604686638, 0.0318717318944651, -0.056816977384796, 
    0.0460870772736808, 0.52414287425662, 0.0188191012823484, 
    -0.0294145704953852, 0.0762997493542794, -0.322156239577889, 
    0.685076983574573, 0.325226668805654, -0.190180933134941, 
    0.535340828670686, 0.449760241049646, -0.189922116884446, 
    -0.149013604389261, -0.305472424785107, 0.767706580808529, 
    0.146165683735975, 0.130811896384639, 0.0550888663846692, 
    0.727468456171245, 0.00351501663330983, -0.0637272432860449, 
    -0.00929986903329523, -0.379054692024717, -0.0851766628304659, 
    0.264947051295071, 0.185178854013533, 0.222617294179651, 
    -0.00984337838209619, -0.350976253429479, -0.415556673279122, 
    -0.000436745610573927, -0.301747006993283, -0.247590362418951, 
    -0.100440108746688, -0.297031970917829, -0.0771688098271535, 
    -0.212572083688168, -0.0360342635644246, -0.250769245194154,
  0.0462825758265188, -0.00686474049911796, 0.0238756595045142, 
    0.0309661407992365, 0.0113714465573383, 0.0391009413964229, 
    0.0422818885771138, 0.0758943195597571, -0.0131990941402512, 
    0.0134050449008437, 0.384805857854694, 0.337546061623757, 
    -0.113682536451797, 0.61730639527437, 0.399083015613049, 
    0.036331388103915, -0.14781090457627, 0.937579878065621, 
    0.269758473741906, 0.0691526612088479, -0.463598084976326, 
    0.0150675966824856, 0.89423214906631, -0.0119698800466003, 
    -0.15865408005613, 0.0771222426258135, 0.943418577047349, 
    -0.0974091598026854, 0.541814424107348, 1.01827188711895, 
    -0.0423086012519358, -0.00172603912774502, -0.0600943905279634, 
    0.000456018147199033, 0.0463611211839686, 0.0196078857360423, 
    0.00934814278849505, 0.00263563018053997, -0.0930856582518479, 
    0.114905408145741, 0.28249689766344, 0.0198937258915567, 
    -0.102908606033601, 0.0615644055320293, 0.422901287564313, 
    0.405397341413002, 0.144627731711137, 0.229258715529628, 
    0.717574308315754, 0.161898717793482, -0.015958777903077, 
    0.0264121796087894, -0.0978300287562149, 0.296968462364408, 
    0.192178617957154, 0.160208833758523, -0.0604925807305422, 
    0.24600887814178, 0.160720703408771, -0.0621694309109033, 
    -0.101738521923665, -0.264172946787559, 0.0854815724240311, 
    -0.226901127526836, -0.0546707959519939, -0.0594251279395536, 
    0.103353982201128, -0.152644969180255, 0.127745505967962, 
    -0.296454847598063, -0.0358049150166129, 0.0356714797530827, 
    0.10112967381109, 0.0775590309984583, 0.0398891602799216, 
    0.0737273499390053, 0.064039305954184, 0.0612505295665307, 
    0.0710065414083442, 0.108870532624015, 0.219111544503412, 
    0.053861936883059, -0.0177935784540015, 0.361530214439496, 
    0.343944822127214, 0.129774766127476, -0.0291288695440742, 
    0.104809408192661, 0.257950713295297, 0.168634458630149, 
    0.363553687841062, 0.522132756749502, 0.237730063311765, 
    -0.0852212087043313, 0.574059275912974, 0.37869254896163, 
    0.108710011664187, -0.168069373230222, 0.564213642559085, 
    0.345539014393914, 0.0572938292654861, -0.0490615036846577, 
    -0.103214231866104, -0.0688246628682628, 0.653778513588351, 
    0.249589250335637, -0.0911743791865643, 0.277934661669991, 
    0.419612710924126, 0.0884279269698896, -0.0617758762313161, 
    -0.0505702341339268, 0.334874385733923, 0.299415868298458, 
    0.123999779471755, 0.0902234120364266, -0.167767151811712, 
    0.203166500626163, -0.138822133194379, -0.329020297416604, 
    -0.207521603727764, -0.203052718690147, -0.1971385988098, 
    -0.207935812495941, -0.209642828038482, -0.073313983427216, 
    -0.231382777894174, 0.0527036002289815, -0.269497929654357, 
    0.00390217911976211, -0.133833121112306, -0.0246207838660419, 
    -0.0431330672293636, 0.00189170683662174, -0.153970273176973, 
    -0.0309184090765446, 0.01342601158911, -0.106149172017245, 
    0.0129567194881995, 0.0395182012364587, 0.167648130862728, 
    -0.00870357877946378, 0.0794593068281296, 0.296631225884932, 
    0.0846598249313383, 0.022810563641012, 0.0203308915462932, 
    -0.087522526442774, 0.379934293290886, 0.238139256390785, 
    -0.29144644126865, 0.318289492421557, 0.595980304108644, 
    0.137499188455527, 0.657075962125705, 0.670547980770853, 
    0.209759086051781, 0.108750748360852, 0.3142669707796, 0.462441998757234, 
    -0.0690597268451379, 0.73180036939352, 0.381686272354998, 
    0.0412457013848234, 0.0331013502048288, 0.201859285941646, 
    -0.397871772251033, 0.55492063055616, 0.471349442387607, 
    -0.0983094115216184, -0.248340012420339, -0.0725943309509703, 
    -0.244517037011591, -0.283789018316475, -0.187739954062273, 
    -0.0616628945425581, -0.205895155055106, -0.0492575750830472, 
    -0.158607758217651, -0.0766360859338434, 0.123635390238457, 
    0.0651846765684741, 0.0420011559985404, 0.0391417893032613, 
    0.043367492504278, 0.0388144046653729, 0.00703202853081973, 
    0.0799901921684465, 0.113085471789095, 0.0961230109210448, 
    0.356308259871226, -0.110366028306729, 0.436069116554991, 
    0.511852022011248, 0.145603754618347, 0.0305608663927376, 
    0.374109356642762, 0.369725384834829, 0.318859420717919, 
    0.268709748972871, 0.060103106919237, 0.345561534953475, 
    0.527932881015785, 0.274188283742193, 0.0773559533264888, 
    -0.0518839663981495, 0.0417957382114419, 0.22958553731406, 
    0.0325609130956851, -0.0774809395201987, -0.0735935793361443, 
    -0.241837360083375, 0.0204430303959828, -0.0661568431493758, 
    0.0541486633770909, -0.104468780363188, 0.0772281499621791, 
    -0.109296836644068, 0.0490704941666426, -0.302441116381535, 
    -0.0142093964430721, 0.015351680825335, 0.105029297045869, 
    0.207224892560108, 0.175124722401198, 0.0797867324144288, 
    0.00116221816337957, 0.106783688813893, 0.226592219937447, 
    0.438675436507833, 0.327402664852288, -0.0721634011865187, 
    0.213670252402436, 0.825572741818094, -0.0722902256898887, 
    -0.129613991374487, -0.0754469145504346, 0.793180581082147, 
    0.213036379860863, 0.26040163972544, -0.26970681686369, 
    0.413875824763623, 0.515521519219014, 0.2723926748016, 0.020610318357077, 
    0.641237512693103, 0.344924483955274, 0.144376367207821, 
    -0.207717036305515, 0.296122597036862, 0.428030459210051, 
    0.301440546640974, 0.205465283998427, 0.0924757841201279, 
    0.294942405903287, 0.547878131944138, -0.29875761764442, 
    -0.324885377726676, 0.102032603334545, 0.313277091762059, 
    -0.0763126307582914, -0.0374212668068098, -0.0142649922339743, 
    0.0210185481537307, 0.0205267625458602, 0.00534951812831036, 
    0.00306054277311124, 0.019301290518282, 0.0250166872475714, 
    -0.0970430026073884, 0.153421693687795, 0.189132419365006, 
    0.0604088253052497, -0.0359321608508271, 0.27120054725556, 
    0.314779301689529, 0.105398775685377, -0.0017557109482496, 
    0.0298146084560729, -0.140820799708493, 0.631239459657844, 
    0.275449830409086, -0.136614019766901, 0.174885120579184, 
    0.554843857851908, 0.245375660619784, 0.124227348793536, 
    0.154549462122538, -0.0829981161280602, 0.318007336074886, 
    0.553180411321022, 0.234579920078427, 0.0622477546955113, 
    0.051259588116812, 0.0614468959993632, 0.0173467443124179, 
    -0.121201922454678, 0.212243349853947, -0.00617818110181578, 
    -0.100114950432139, -0.0062070973785496, -0.194533536047845, 
    0.128151915419639, -0.212407722942207, 0.0300852836252825, 
    -0.211382789173443, -0.0133867305723315, -0.0798536570682705, 
    0.0792554352247095, -0.310502062116216, 0.00718159471536528, 
    0.0693502978456741, 0.0821684037740635, 0.0932158020567446, 
    0.140709140194955, 0.167668133348416, 0.195194847421651, 
    0.260701985410352, 0.186441817947452, 0.0489906003817119, 
    0.00258905080988364, 0.24450953104292, 0.457800715845782, 
    0.38720273216676, 0.28870841951006, 0.185584213465735, 
    -0.0520743556813969, 0.430942425704799, 0.86521706405665, 
    0.173847214740804, -0.264222054028559, 0.213682111203094, 
    0.386231039460667, 0.364145996085786, 0.68860997807068, 
    0.0302777277122308, -0.157094777980772, -0.293101443885513, 
    0.131962288361849, 0.415598803650421, -0.236367871700389, 
    -0.0531807284136296, -0.0828579156556754, -0.0844325074095954, 
    -0.0722777078632103, -0.0849117832133446, -0.0826753153944165, 
    -0.0790875534687004, -0.0515958125232382, -0.102313424534481, 
    0.0420271033673965, 0.0513620267450532, 0.0771893611391731, 
    0.0643495799887138, 0.078199323893217, 0.046082686793909, 
    0.0599266350835439, 0.0672071892643936, 0.0774802196561115, 
    0.0479760836067096,
  0.130059099345308, 0.142567512050403, 0.148046688226242, 0.193890209658699, 
    0.207203682908075, 0.139920165847558, 0.149303211538782, 
    0.297131783424437, 0.186473269591501, 0.0200050870565697, 
    0.096483711390584, 0.291640050074078, 0.202128614357409, 
    0.333897897659617, 0.432936245234913, 0.147200585479365, 
    -0.0958579302465895, 0.393267914261608, 0.48351656149456, 
    0.313785833853791, 0.270632805423628, 0.271443186940496, 
    0.170470902101412, -0.0304281318423071, -0.0189927624086884, 
    0.482261225326896, 0.773376878889004, -0.345965585980263, 
    -0.345939960569343, -0.00817102655545891, -0.256932094862433, 
    -0.180400649420376, -0.203209186241588, -0.236496276864154, 
    -0.144742783261397, -0.228437204214278, -0.151078458968456, 
    -0.179810334397925, -0.130947646510019, -0.135738550864199, 
    -0.0280529687819735, 0.123892924981263, 0.0538484483147607, 
    0.0784977481544703, 0.0734093440118761, 0.0935994569922423, 
    0.0805190817941803, 0.0735391764221651, -0.00800835222116503, 
    0.0199674334065363, 0.0819892167946937, 0.0867226998995147, 
    0.0902195524793523, 0.173516574160616, 0.139986124082247, 
    0.0389438543818168, 0.169246903560284, 0.213951765054448, 
    0.00378843709483731, -0.00652049594841644, 0.404176796285595, 
    -0.0581737678888277, 0.64314662773802, 0.346527904767481, 
    0.0691675602116728, -0.187759006308034, 0.494911870310748, 
    0.46026899060647, 0.14673032024069, -0.0771015736550501, 
    0.127967295437256, 0.472438681056775, -0.0988762266256403, 
    -0.0363166918411793, -0.113932193363837, 0.363693979076351, 
    0.0742839130362439, -0.107211509640078, 0.228191293896151, 
    0.178753079970347, -0.135655779968863, 0.011059015386677, 
    -0.217593400937306, -0.0370868584295903, -0.192927782312381, 
    -0.140066203973858, -0.0443772619201008, -0.0388852616474392, 
    0.0104808847082996, -0.160563390683383, -0.136042268927158, 
    0.262612089914683, 0.147001791264299, 0.0461819200845386, 
    0.0308576746543799, -0.207979796145445, 0.342751016472205, 
    0.356352528656726, -0.060212257893685, -0.262805080346828, 
    0.0472178405887074, 0.466709542924344, -0.0621567387878086, 
    -0.284577323965941, -0.164045013538139, 1.1743235680193, 
    0.37895560753874, -0.0579978536172276, 0.796565880169698, 
    0.129909817151033, -0.316734048839129, -0.166899609240106, 
    0.101985215538635, -0.143043302643585, 0.0998230289408551, 
    0.0729179708106541, -0.0236530274855041, -0.0399233839298879, 
    0.00376444513185777, 0.125121444383952, -0.133266610365654, 
    -0.070439621941213, -0.0318037761505398, -0.027383702433598, 
    -0.132922061395907, -0.0197293512533046, -0.0892826232987125, 
    -0.00694317282510247, -0.0685374392182767, -0.0765548665935518, 
    -0.000110871508559748, -0.140196860344776, -0.00696033449926431, 
    -0.0370221721056647, 0.0344109157760389, -0.0697691524919508, 
    0.0581849531138157, -0.112576298829056, 0.0169183008270858, 
    -0.152078791082678, -0.0259660056169374, 0.0407492337423053, 
    0.0617619737578484, 0.133102141533127, 0.177092747475059, 
    0.0763220206830308, -0.0558219963368346, 0.0579721689815746, 
    0.369151560663903, 0.0602457089967755, -0.0185629381713339, 
    -0.164449856250241, 0.678813216732956, 0.277525283875906, 
    0.0921384694669397, -0.272659263662412, 0.139405156807973, 
    0.60231982570793, 0.224375090407253, -0.127616240405952, 
    0.528089146490474, 0.582576811147627, 0.0929648897590124, 
    -0.0603470457605335, -0.1503676680246, 0.537328456464434, 
    0.248977924832215, 0.00159799553272677, 0.539489524152512, 
    -0.0981914927792382, -0.441828169893671, -0.132669217174653, 
    -0.123991722165616, -0.184048572454266, -0.135722616243277, 
    -0.0954727112809982, -0.06134672659397, -0.135045449641212, 
    -0.0357221998080521, -0.188981830516673, -0.0816980066652065, 
    -0.0622686213220607, -0.308380618310508, -0.140670165524245, 
    0.085021781876034, -0.173813021861798, 0.0714278339335252, 
    -0.046932335162632, 0.0401699424658904, -0.189558782544033, 
    -0.0133289011962637, 0.0555850334475483, 0.0709234670266268, 
    0.0542032553492582, 0.0589296682566223, 0.0525075562044123, 
    0.0569640909707355, 0.0622244384904423, 0.0606140874481361, 
    0.0422483743724336, 0.112239174279389, 0.118854868638795, 
    0.113047137423445, 0.122213645844755, 0.128220537273685, 
    0.110468576329526, 0.110221131618079, 0.144744401393335, 
    0.135082683085106, 0.0824602120839522, 0.0782955653347365, 
    0.154016751213472, 0.280131358892771, 0.158562096511409, 
    0.09558923037568, 0.440371986368568, 0.279076893679454, 
    0.0537260975576382, -0.182331345502754, 0.103285087762501, 
    0.560925622133001, 0.18627767647112, 0.0335146528756636, 
    -0.193018154627517, 0.274094407390691, 0.535449824704208, 
    -0.165151162161216, 0.625111800684878, 0.782755815120685, 
    -0.090282833617156, -0.120605611877885, -0.280728073881441, 
    0.0145869390595073, -0.0892941017724617, -0.105311192521305, 
    -0.19399560628378, -0.0449540131949155, -0.149999399268609, 
    -0.153427117175795, -0.0978597503930769, 0.0934667566506253, 
    -0.231649727256744, 0.0557594701879854, -0.135161653215546, 
    -0.0452158044637321, 0.00939543138235978, 0.123725758510366, 
    -0.136343202291078, 0.044879146429771, -0.382337456235919, 
    -0.147942780290138, -0.0340842336660302, -0.0968545384172908, 
    -0.0497402166846557, -0.0033077030535327, -0.0859967363336831, 
    -0.0031335885765882, 0.0401786365681015, -0.0557418487684649, 
    -0.0362264796158221, 0.158521644113685, 0.329088655674536, 
    0.103151787415286, 0.866622094807219, 0.0915126909574286, 
    -0.0768028948545655, 0.041470488152525, 0.220937115538109, 
    0.29198136196586, 1.04844451068881, 0.296233080766212, 
    -0.059346370829744, -0.0518350818963579, -0.012061871461385, 
    -0.0864905128845392, 0.0332152366507921, -0.0410967547082552, 
    -0.136619902644346, 0.0213539089979785, 0.0235839212082983, 
    -0.0879035881164436, 0.0543771280228893, -0.0839889191000889, 
    0.00377379180736116, -0.0705593742685945, 0.0169570915943882, 
    -0.235975948114841, -0.00483593041350838, -0.238973650235341, 
    -0.155871338473797, -0.0197285070900724, 0.0596867937536123, 
    0.100837570310097, 0.100541877525403, 0.098334678271725, 
    0.0975170761858208, 0.111369667793011, 0.136250993107792, 
    0.122799377354376, 0.0873632676502658, 0.141019258272986, 
    0.165044804941492, 0.181751515236162, 0.209852715571165, 
    0.199485295371639, 0.149254990616846, 0.201280873424398, 
    0.323915039420671, 0.147798255456611, -0.134013431442494, 
    0.073823101410117, 0.520752354445001, 0.2416989965003, 
    0.0376191933982813, 0.111831437727456, 0.469074587186134, 
    0.131473660101212, -0.13641051014532, -0.0817308291910082, 
    0.782705145554546, 0.296819476772878, 0.0104589016413613, 
    0.255293489663236, 0.519969333857561, -0.136517380669709, 
    0.454654709925798, 0.508377052094695, 0.605622742632656, 
    0.925081578183587, -0.0252172550703881, -0.361399018811115, 
    -0.13317838403519, -0.0804457238191438, -0.216108378473493, 
    -0.0970640880309669, -0.18111265610484, -0.191287813535946, 
    -0.133242097924798, -0.0410783439710789, -0.243777253025042, 
    0.0825156739212749, 0.022768496675956, 0.0611883707630204, 
    0.0191933696536334, 0.0562893459279872, 0.0143330002705953, 
    0.0682952691599194, 0.00937925697128349, 0.0793068578799812, 
    0.000961459876834145, 0.0563621611313685, 0.0961517986569547, 
    0.113341136518338, 0.115576514544255, 0.117795522562902, 
    0.115205525732232, 0.113983922964099, 0.124553785578098, 
    0.117982109984602, 0.0950497115341044,
  0.0295863217883575, 0.0602568144871337, -0.00173646154617016, 
    0.0756325314144654, 0.187734154084186, 0.108407615715597, 
    0.0672995174693985, 0.0718891931106424, -0.0494651452849252, 
    -0.115857153929536, 0.643176928311356, 0.184133528407058, 
    -0.0795323930860599, 0.22976777259965, 0.154145235468494, 
    0.0493135388155228, 0.948683554600273, 0.450418283173539, 
    0.0479146613572037, -0.248647339348944, 0.0580358127192388, 
    0.871779754610431, 0.0663766854384268, -0.211904492898367, 
    -0.257673251316387, 0.377785478635521, 0.592454162304411, 
    0.241300846116069, 0.0104884225713004, 0.0131086035510986, 
    0.199712311644469, 0.181348278372641, -0.173721928257527, 
    -0.13993826040584, -0.104761358415876, -0.0693467109804736, 
    -0.0290203599653838, 0.00985483244477343, -0.0664739316849818, 
    -0.131125076490158, 0.160361191517228, 0.0907563348316138, 
    0.0455516298330007, 0.0369643647754105, 0.0474627488125044, 
    0.0545417510724908, 0.015110177822536, 0.119173422316291, 
    0.0219486556796746, -0.0247967241551107, 0.259364863183648, 
    -0.0277452083497608, 0.500331934086694, 0.298634244339823, 
    0.123967822896768, -0.104005353377629, 0.461300656024198, 
    0.278749949703414, 0.0105708648657619, 0.375185131485661, 
    0.382550416129902, -0.0127576379174785, 0.0300890165841798, 
    0.0048029132056084, 0.292557354747172, 0.127135529124111, 
    0.586465043818935, 0.250313269731691, -0.106997468292884, 
    -0.0828184188196314, -0.219022502181627, -0.264735323664803, 
    0.0498397977622699, -0.0661742072885812, 0.104134449406981, 
    -0.200669155519835, 0.0666639411450321, -0.16381778039132, 
    0.0835053260041963, -0.278119111779325, 0.0221440592943523, 
    0.0822842423982546, 0.173273633413921, 0.179562320827423, 
    0.0888856615374611, 0.149448931014372, 0.405399724611066, 
    0.373074804973159, 0.191270501242565, 0.0720833895639778, 
    0.2133267867061, 0.41841756296561, 0.373052984955077, 0.264813921993864, 
    0.298289463927273, 0.468697760968343, 0.475570173242061, 
    0.250515073596989, 0.0101733648504435, 0.181750979288983, 
    0.625409522310218, 0.270636019860024, -0.00250483366596109, 
    0.374193686808817, 0.370168049903215, 0.0977845070160605, 
    0.378949437732363, 0.551963086514307, 0.166063326995771, 
    -0.197588348952897, 0.466186517953004, 0.329665250197735, 
    -0.00479253159557663, 0.0740418448935567, 0.654057861789583, 
    0.439941257919646, 0.0506401409609265, -0.0175675647702087, 
    0.106925364310579, 0.674060064329604, -0.362360343829421, 
    -0.13488138489687, -0.157190600782231, -0.205345213560397, 
    -0.128941911808331, -0.191014870882057, -0.137003283563238, 
    -0.113048990192432, -0.209145894587378, -0.0716643757240738, 
    -0.0245826931083469, 0.118584485927318, 0.0407489956179253, 
    0.101373372094732, 0.0294173503587632, 0.101360311395668, 
    -0.00465673053725413, 0.0773414194921293, -0.033815333165061, 
    0.0293872134940626, 0.00838961232306314, 0.0384404124730572, 
    0.0159662238148267, 0.0236269817763947, 0.0701078087833516, 
    0.0107880133067056, 0.0384550895159576, 0.0471560498558998, 
    0.0544953930352895, -0.0132214971641791, 0.0541684674795372, 
    0.1261216261119, 0.123153589597875, 0.100846916872294, 0.133905415740611, 
    0.205442463225711, 0.238046544134761, 0.131020065354744, 
    -0.0176381706332878, -0.02347453984279, 0.497696851241291, 
    0.246006975865327, 0.107416632465949, -0.222128611745918, 
    0.133935050340648, 0.598219451029175, 0.302068687956483, 
    -0.125641812765029, 0.421790348112832, 0.375789871785238, 
    0.0592632659048271, 0.0278530970004334, -0.0571801799850997, 
    0.582805049646525, 0.0394049238134183, -0.309317672653541, 
    0.140322400159099, 0.491679831270963, -0.0943795005874995, 
    0.0375601089887248, -0.344166475318124, -0.0402294858977454, 
    -0.238347700163226, 0.0630891081996829, -0.196571925828041, 
    0.119612407623787, -0.302051861852043, -0.0141027666492728, 
    -0.267550022672202, -0.193521984365435, 0.00362488639713032, 
    0.0766765956040775, 0.0419062920520152, 0.0747847534130917, 
    -0.0428292410185785, 0.0258421522893503, 0.0281223836192893, 
    0.066900384576696, 0.0622169946178028, -0.0138682395361942, 
    0.0435654546725065, 0.0760942120374976, 0.0859519519439787, 
    0.114830384429045, 0.12815832135931, 0.103522368219781, 
    0.110144599414681, 0.156025025188509, 0.102739869646861, 
    -0.0098573000973838, 0.36530884167833, 0.206495537680423, 
    -0.00785413032729738, -0.100026086799414, 0.372157974541849, 
    0.367879074054116, 0.226079704222066, 0.168199555840219, 
    0.0895534757974114, -0.213976941374533, 0.0503498934348839, 
    0.59491401192117, 0.282062195097076, 0.043342274030641, 
    -0.0147298518463704, 0.310571701602921, 1.02953223712606, 
    0.0128106515651765, -0.368007085266081, 0.0885142209996514, 
    -0.313450713393133, 0.131964559976451, -0.323921558140054, 
    0.0611707238923585, -0.35007739916117, 0.00188987361961561, 
    -0.333184746318175, -0.098297509163555, -0.211615098006264, 
    -0.131971741235617, -0.0552939714013595, 0.116008535959898, 
    -0.0734577964169627, 0.047140501021558, -0.0150392976111581, 
    0.0499692082066043, -0.106462956783917, 0.00712234634406508, 
    -0.109960330134276, -0.114998556105775, 0.0416416395895494, 
    0.0484083598402134, 0.0618170638782521, 0.098705556169866, 
    0.117554709828482, 0.103742060415771, 0.104059876628618, 
    0.143412397798002, 0.107225792806118, 0.0383566490939721, 
    0.179009818859269, 0.153935822153625, 0.0494287346497743, 
    0.462367963306263, 0.355445120924306, 0.0331911870737005, 
    0.025098881324439, 0.591745320577531, 0.349359208671391, 
    0.180329084315776, -0.259383984004596, 0.353258993658676, 
    0.46890404474363, 0.120133590690475, -0.0151120385446737, 
    -0.140956222250955, 0.0435409821381297, 0.376801582036175, 
    0.635005758859421, 0.297549738892727, -0.107945371484903, 
    0.345452023455689, 0.337161016279248, 0.0302652743110856, 
    0.0326734584982742, -0.217614344045605, 0.334501057028287, 
    0.22286919644552, 0.109063142760856, 0.299230314901494, 
    0.088725437004853, -0.0314054451355556, -0.0552598499777237, 
    0.0931803416737556, -0.0960962983292232, -0.096435459288739, 
    -0.0276840252682619, -0.0749639571139602, -0.166429345328013, 
    -0.0651927030093424, -0.0951840985249707, -0.102182174237835, 
    0.0845101034324508, -0.103184551860276, 0.0397989989145673, 
    -0.0625804039795021, 0.00772769871619941, -0.0395050070360065, 
    0.0337429844742246, -0.140712051753827, 0.0116640827179719, 
    0.0732059232687974, 0.0807669506555616, 0.129581960388174, 
    0.148227937801812, 0.06461466778851, 0.161644722840955, 
    0.303843978136386, 0.119085193410846, 0.095114501362864, 
    -0.199494937647667, 0.406754423806916, 0.349393278712486, 
    0.166463799860142, 0.107485754298234, 0.0223311706616319, 
    -0.190874370392671, 0.275989694368726, 0.673391208486931, 
    0.455855264035276, -0.0027320570709721, -0.216398981089468, 
    -0.297495697657165, 0.203994390931267, 0.52925005855091, 
    0.263338708339086, 0.0160463396396663, 0.612255505550519, 
    0.227660695901226, -0.0503914958344181, -0.191453399560789, 
    -0.000525699955527523, -0.130680838343527, -0.0496901426859175, 
    -0.149494660864084, -0.127230305115544, -0.0987423953551242, 
    -0.16536755373493, -0.113020049005431, -0.0822041718760934, 
    -0.16902420586693, -0.0107761165157575, -0.0830818598303918, 
    0.00531743693599845, -0.203863627958555, -0.0638568796357585, 
    0.0251221778884939, -0.0316424952093168, 0.194297509531763, 
    -0.150876931637938,
  0.0399823634119584, -0.0220423184618187, 0.0474354793818918, 
    0.00711434247380455, 0.076024772907839, -0.00710201697470153, 
    0.0471522941683753, 0.0289054736416733, 0.0625948285976368, 
    -0.0361569153970674, 0.0434523668938361, 0.0770720488800982, 
    0.0911892332847754, 0.104910999491378, 0.104420333689303, 
    0.0908048689339809, 0.103650797148037, 0.166762992086315, 
    0.141666630119643, -0.160132092047, 0.288497071892422, 0.303575078455791, 
    0.0519960843079991, 0.351042536704534, 0.359338795135105, 
    0.0521448092673549, 0.382755739014424, 0.593781668419493, 
    0.180120167561013, -0.268263962872259, 0.449141377288487, 
    0.498238125336304, 0.170567311578464, -0.201009409540817, 
    0.420763661296662, 0.399739237313155, 0.193459135315316, 
    0.565842613492946, 0.370331578582548, -0.0142449775807851, 
    -0.161546867143526, 0.0621126200465651, -0.122595751950868, 
    0.0375189831769453, -0.28936904768917, -0.0844914743762706, 
    -0.0405247740078033, -0.146318728395937, 0.095807114824419, 
    -0.195944247743701, 0.0169198049549199, 0.0797042222853403, 
    0.136644869186687, 0.236352413552877, 0.249990590368505, 
    0.189724695582186, 0.18678406861635, 0.276202665377062, 
    0.293019666185411, 0.250810488616636, 0.271457933699587, 
    0.308078059689975, 0.315635038323108, 0.261787617900866, 
    0.199071823007337, 0.318716683056564, 0.469735838730069, 
    0.264629963782914, 0.00249733696535881, 0.284946754214554, 
    0.56669223868363, 0.206959409068711, 0.0388292231131278, 
    -0.178785480568529, 0.0151761768112012, 0.689486354694829, 
    0.300027920868425, 0.00575964325413649, 0.603783440705941, 
    0.161889992024693, -0.199625948370221, 0.191042311410387, 
    0.495274831836605, -0.351996738633306, -0.354945557989332, 
    -0.0305210797001393, 0.0418259894268767, 0.518506235427389, 
    0.624411594650985, -0.183997321344664, -0.307363131840062, 
    -0.106099178473576, -0.134123207742422, -0.182274493176607, 
    -0.118725390889961, -0.102275333468543, -0.132914419324297, 
    -0.11523498195308, -0.0739682425838721, -0.178107853424161, 
    0.0488675108565416, 0.0269344013805206, 0.0603935193895864, 
    -0.0123748310327673, 0.0331677316175098, 0.000758340843766706, 
    0.00286962689905484, 0.0376029480791297, 0.0766732761362168, 
    -0.0850355403641837, 0.126864725819009, 0.26619440147701, 
    0.163923488248958, -0.0878764943417799, 0.380638806518433, 
    0.40372965115627, 0.131902982951966, -0.179058915102163, 
    0.413761781123226, 0.297699391917502, -0.195748277744004, 
    0.0325293110178499, -0.249978643372302, 1.10378629642014, 
    0.60097668009441, -0.562312437136335, -0.196951650442224, 
    -0.515106028524902, -0.00294616930542788, 0.617946347533294, 
    -0.352216931432433, -0.0711559961294622, -0.05400925092122, 
    -0.101404151830311, -0.0497427762687133, -0.0427200040677452, 
    -0.0602644078347157, -0.100748413923085, -0.00965800802596706, 
    -0.0969627110286024, 0.0694551962033464, 0.143211782572533, 
    0.122339397072802, 0.104697949107416, 0.115015564260636, 
    0.192068491976885, 0.194585084142839, 0.12921401831846, 
    0.0919057935776477, 0.121780990127533, 0.162711012959547, 
    0.16169693586961, 0.152930806992454, 0.158240682778605, 
    0.163166534922676, 0.145788921395616, 0.118739129867462, 
    0.163437169756569, 0.239493432568297, 0.198376226398722, 
    0.114763202738426, 0.0889651543655368, 0.0992163683406505, 
    0.115782225972591, 0.129935583668105, 0.107232540662795, 
    0.100178780149742, 0.13830051911248, 0.122309246168371, 
    0.0826787632084401, 0.158633526509684, 0.127840918755513, 
    0.0759910594115721, 0.354119198442251, 0.273077191342416, 
    0.0380994431256285, 0.0308629782476172, 0.429478715267867, 
    0.310106379841785, 0.0825620542014049, -0.0756590411766301, 
    -0.172770087657171, 0.338454539423111, 0.391813546664936, 
    0.33558568116726, 0.152627347047271, -0.103928700948134, 
    -0.224127548068174, 0.314780124768719, 0.569252423523456, 
    0.209377242736831, 0.0239299413501731, -0.0712486844663872, 
    0.421415132204973, 0.288062723431807, 0.0925709494269032, 
    0.0642403754645476, 0.154037058401209, -0.161338706351383, 
    -0.190339486966914, -0.208275118869401, -0.21113821201222, 
    -0.208630198598508, -0.190419880225904, -0.150978283958241, 
    -0.19927978064944, 0.00142514236799163, -0.193094443938892, 
    0.102658294565736, -0.204712402019157, 0.0622905994606534, 
    0.0122801208073476, 0.0429566763882175, 0.0459554584736566, 
    0.0651860039367203, -0.000173154399672359, 0.0516778825387532, 
    0.0378483787988539, 0.0577534904040453, -0.0398900513066959, 
    0.0465793150004887, 0.109195229924724, 0.0710462792444468, 
    0.0980846540773326, 0.226996626878715, 0.141349041564356, 
    0.0100827472429456, 0.0658922170267588, 0.27302847225952, 
    0.237160774172206, 0.214588277908016, -0.186101607734377, 
    0.165590305241179, 0.499065182493077, 0.242118396059386, 
    0.235876013859721, 0.298883048051864, -0.318607540924487, 
    0.29382059974809, 0.498450198961982, -0.214478241417732, 
    -0.270410021527416, 0.00932593380220458, 0.238598899185598, 
    0.0930650614551308, 0.0952875014103217, 0.158362777364841, 
    -0.255621226490091, 0.220684445955471, 0.148715131452576, 
    -0.103143958951116, -0.00105168317509349, -0.187585992071921, 
    -0.00143571844703823, -0.326138066178798, -0.104621657053257, 
    -0.313174000017288, -0.298074821537648, 0.254427947394043, 
    -0.25754621361057, 0.16313858235637, 0.00782386389326875, 
    0.0267452289220262, 0.0493111028718662, 0.0794207884483915, 
    0.0592659279916779, 0.0912654206508407, 0.0786641158565603, 
    0.0678122202351584, -0.00309038316066622, 0.0527233142409539, 
    0.0927707618490625, 0.0934396306511399, 0.1288345711411, 
    0.185535898280761, 0.150135067248449, 0.120145444574347, 
    0.119147690305688, -0.0221389248811296, 0.14071188824621, 
    0.481766711979878, 0.199927611964955, 0.06949179894099, 
    -0.0017478514786619, 0.0378396862355013, 0.282284926922138, 
    0.00118471322652182, 0.4925461824332, 0.920909492631605, 
    0.0915526192369726, -0.307296058751225, 0.149667720048819, 
    0.314916197654477, 0.289480944526716, 0.549373471330623, 
    0.216513319667177, -0.00580369578184807, -0.250627044948931, 
    0.274035958074444, 0.0274966719961395, -0.216823366867333, 
    0.086700140028587, -0.340418567510399, -0.0442415835690143, 
    -0.298656074378716, -0.240355561986292, 0.0839188882279669, 
    -0.247648514433547, 0.140693624038937, -0.22279615499581, 
    0.0928359975624961, 0.0145352767222262, 0.0676367981012588, 
    0.0117939938315745, 0.0536441154458931, -0.0304032916320704, 
    0.0281596932575154, 0.0272110285054002, 0.0409175000310848, 
    -0.0609769465386403, 0.00952547551998553, 0.181498651719207, 
    0.060739389375574, 0.0363876784367047, 0.311413789693106, 
    0.148735443798469, 0.082105341669299, 0.208374247157791, 
    -0.136366865657006, 0.393174252650977, 0.486859296265545, 
    0.0930369032478068, -0.190050267896228, 0.848472729572824, 
    0.241728074218378, 0.0924456208040789, -0.241283631897749, 
    0.208837599397112, 0.410721417818338, 0.466926823057309, 
    0.543957666689956, 0.306352504717268, 0.0493268352593593, 
    -0.00739505049595538, -0.0144217429676503, -0.0181242108499599, 
    0.223472062144403, 0.375217835525016, -0.128320746135393, 
    -0.152500743155236, -0.144254906548233, -0.210006721910473, 
    -0.12211556421141, -0.234790242313826, -0.150479868063321, 
    -0.238112024992951, -0.0889078546044994, -0.254580080788811, 
    0.00304000654245687, -0.202092727900066,
  -0.16781933605864, -0.032118005673358, 0.432824989064039, 
    0.245049310517991, 0.10035380000325, -0.217090554582517, 
    0.023957386143998, 0.440898193757555, 0.128370707095787, 
    0.0305401501267392, 0.0728450012594697, -0.23594016697028, 
    0.198694123500207, 0.515824930421224, 0.214975457409866, 
    0.164611143292833, 0.282157967312513, 0.26921387003302, 
    0.529540732440538, -0.210181053770436, -0.333382532403972, 
    -0.0398390446391212, -0.26931420204371, 0.0105958893863611, 
    -0.296970852073952, 0.00448180852123893, -0.328562928466393, 
    -0.140259641386571, -0.104023389499667, -0.270428620257102, 
    0.0413030258487579, 0.0908100095011364, 0.0958285359175292, 
    0.0930123713535765, 0.102964607696542, 0.0982725309785483, 
    0.121929821958321, 0.112685918640447, 0.151301698258075, 
    0.134483073211567, 0.0940165848477144, 0.0623840751324246, 
    0.0706226251402638, 0.0767773696801371, 0.0841265685314902, 
    0.0553731001679497, 0.0710199243073966, 0.0864229503115565, 
    0.08680152387088, 0.0241247330991202, 0.0584948779228725, 
    0.138772658380902, 0.173659431367529, 0.144693485229684, 
    0.0948142608389627, 0.134131162155023, 0.255135394366074, 
    0.220511218441483, 0.330159549885639, 0.267978355211318, 
    -0.213006499252394, 0.264351502547727, 0.50867016248963, 
    0.202889921392309, 0.118843792950651, -0.279269280439617, 
    0.324946737226053, 0.38946453688465, 0.23259794879799, 0.476271425872815, 
    0.322030062908575, 0.133660090476996, 0.0635603168227293, 
    -0.0470974235793511, 0.223565710555987, 0.0206832000185684, 
    -0.179075311158191, 0.0460502040944431, 0.189295339818272, 
    0.00552881360289498, -0.0687945414834806, 0.00544342958509035, 
    -0.295757814729442, -0.0730136629280773, -0.198959466563737, 
    -0.31542810767748, 0.189261899340565, -0.104638041174908, 
    0.121815442804226, -0.269624879903459, -0.00910204771744377, 
    0.0352108750586936, 0.049236577886903, 0.0713265799985606, 
    0.0835446091342229, 0.0686606108852796, 0.00257297218841648, 
    0.0407040729748766, 0.0553743529861782, -0.0110917931876357, 
    0.124222214932153, 0.149083422491555, 0.147737305194666, 
    0.251457531297641, 0.196631667048296, -0.0219135198377267, 
    0.347740478422488, 0.322201821881302, -0.151130710945128, 
    -0.146070193116978, 0.467641045194218, -0.403906096617924, 
    0.35931756908587, 0.477719575474089, 0.469916045637943, 
    0.944527101973339, 0.345588914136907, -0.106806986306257, 
    0.547045292227677, 0.548644981632615, -0.347740607808247, 
    -0.124752860812023, -0.148410848168052, -0.134276153152077, 
    -0.198783876671467, 0.0348627765449687, -0.0181145294868027, 
    -0.0696353778184687, -0.114561351398306, -0.0511518585381054, 
    0.0364986575582167, -0.021627355214853, -0.595487929252236, 
    -0.0408480560301599, -0.0301709474964326, -0.263068954390593, 
    0.244483092001223, -0.168718580755893, 0.12882641606124, 
    -0.29213096358253, -0.042566049352538, -0.00868840731006994, 
    -0.00232208660766676, -0.000956521856277537, 0.00449682558049257, 
    -0.0025508525033848, 0.00489818566966031, 0.0586057581416844, 
    -0.00449114259334629, -0.0431310503624371, 0.458976920444206, 
    -0.0632839495986839, 0.360509456848559, 0.557769015705026, 
    0.185820825537494, -0.0775249352565699, 0.337394511184836, 
    0.271168918737161, 0.0441681898238911, 0.751923276640793, 
    0.480059690110275, 0.0778349866893185, 0.15465501958248, 
    0.675652140868507, 0.154353144831661, -0.153806006147175, 
    0.159517167896203, 0.432444476453803, 0.257433951660534, 
    0.238492346341208, 0.300411388421023, 0.235676525525945, 
    0.12827840699985, 0.0885866766522166, 0.0731639813166928, 
    0.0487724857088918, 0.0540519511010423, 0.131735598492029, 
    0.0826425949477238, -0.136697713255395, 0.132376905261098, 
    0.345683126676724, 0.102348320288106, 0.00160132220394434, 
    0.132995799170284, -0.195529744310436, 0.220980417365449, 
    0.690417701180596, 0.118579220450345, -0.134098821323613, 
    0.192886353730858, 0.317817292649084, 0.0768840094649341, 
    -0.035797515780181, 0.318422897263711, 0.216761867473368, 
    0.239790742876635, 0.394094492585248, 0.160459142920073, 
    -0.0212596042156895, -0.252723394394809, -0.0399739495482248, 
    -0.155640397077067, -0.186776983003953, 0.151672982620192, 
    -0.24486166659821, 0.0054625109676808, -0.118604674401402, 
    -0.0190107950592369, -0.194939084849963, -0.0618683088404524, 
    0.132786731242066, 0.164568840101021, 0.11667938515637, 
    0.121580753898955, 0.0783202045222256, 0.199668216306549, 
    0.445842064847926, 0.32120442058121, 0.141315440774502, 
    -0.213520453077782, 0.444142559229162, 0.488649036291114, 
    0.186398999801367, -0.151948004011396, 0.69844103069402, 
    0.288778770910849, -0.105815740823273, 0.301494296639714, 
    0.54677581802077, 0.116738643976221, 0.195225958001627, 
    0.595933628023139, 0.180815047438087, 0.136987613133896, 
    -0.191052314057171, 0.513585491274257, 0.237329549349682, 
    0.0488124542406534, 0.0201835782765087, 0.205156550666859, 
    0.295992070514394, 0.0705819940812576, -0.0385396076940296, 
    0.0467275978674355, 0.0194572521650416, 0.0287455595660958, 
    0.192733591921346, 0.267254113487251, 0.112529073895489, 
    -0.0267776089861538, 0.00412790038725597, -0.223428262076728, 
    -0.0566486032735715, -0.270717550468586, -0.244683525426291, 
    0.0872046353407154, -0.077161238912084, 0.145511816721113, 
    -0.168936433634727, 0.0761292959882196, 0.0692878336325694, 
    0.0641887962978719, 0.0831000424910211, 0.0915918876572147, 
    0.0793383175634176, 0.0920201359091366, 0.098731233141656, 
    0.0824058498910826, 0.0380427092707273, 0.111279266178151, 
    0.13028864788111, 0.0947339874142236, 0.183992433809085, 
    0.314599040377636, 0.171351191653381, -0.0122245193724501, 
    0.176100797386569, 0.350418394099565, 0.172186135762428, 
    0.259012149588167, 0.26712333133428, -0.261384010491846, 
    0.292844256442784, 0.490644826736262, 0.0649807761814194, 
    0.528324222888309, 0.608826225485155, -0.196043252312108, 
    -0.139005395126584, -0.251927557986829, 0.482785969562307, 
    0.140795674863368, 0.0492603982738546, -0.0445856970729472, 
    -0.0538936063700624, 0.303672011028715, 0.187997539472088, 
    -0.476990900188624, -0.24804008699951, -0.260225767565237, 
    -0.225565472750778, -0.202546446114395, -0.0838858023910247, 
    -0.253555639110704, 0.0572668102066752, -0.115665619284507, 
    0.0691568552712508, -0.354596603592529, -0.0704427610014773, 
    -0.0425793592835894, -0.0974316222275094, 0.0899542622962798, 
    0.0235126643605552, 0.0996107884473034, 0.00464681924579481, 
    0.0547361042239634, 0.042624083307598, 0.0347725575591216, 
    -0.0766811357106414, 0.0182984132935618, 0.0409672223215615, 
    0.056509991672374, 0.0753279019945114, 0.094691139024386, 
    0.0693928550989461, 0.0429562037595451, 0.156266922914447, 
    0.0593792228050365, 0.0806006305469947, 0.340978566575645, 
    -0.184443650247652, 0.247064870421496, 0.487163157987925, 
    0.132519962302046, 0.0847035380195119, 0.153067203342203, 
    0.0103136112233483, -0.342276425456116, 0.340703931491518, 
    0.492640895842633, 0.482774526960033, 0.414920832009561, 
    0.0281297417496583, -0.00603841348219081, 0.958100169609393, 
    0.533553050601055, 0.240619295591653, -0.253468535813998, 
    0.473097322898492, 0.370603565490393, 0.144300995131032, 
    0.0902169871966513, 0.121053612505412, 0.1372656982796, 
    0.0772157272917324, 0.0779740414445892, 0.220719049340063, 
    0.0993065823269419, 0.028689932225924,
  0.1251701264841, -0.0203851006074072, 0.0450703379906573, 
    0.319249836601939, 0.206013764283714, 0.184287934094059, 
    0.267649432764387, -0.146335567657304, 0.410231557999975, 
    0.419276033560122, -0.0798536742930664, 0.41577842813088, 
    0.792886373220928, 0.243058615635451, -0.159199262351108, 
    0.80723955760791, 0.462154135095441, 0.0728988941126347, 
    0.468335226117088, 0.658580444229771, -0.159923190200027, 
    -0.0856007214733482, -0.195105012452079, 0.108056856372418, 
    0.415019759125552, 0.455734639454841, 0.13071864762178, 
    -0.117048987667742, 0.0178539422625311, 0.326989043061299, 
    0.101917848358535, 0.0956297896007213, 0.193563611780723, 
    0.12151493025236, 0.0261661739517178, -0.0384234813913999, 
    0.0612710288338606, 0.042077717650466, -0.11644949784363, 
    0.0662654321753703, 0.191845777058424, 0.0992994830853296, 
    0.0532836264546192, 0.0358195781509543, 0.0449024709582737, 
    0.020016180301366, 0.109359720268819, 0.070151964444602, 
    0.0489138550085993, 0.0362593099784684, 0.00381238159760062, 
    -0.0447630510115877, 0.0328716557479932, 0.0043208914352687, 
    0.0380808239175379, -0.0230200728764853, 0.0381438779487148, 
    0.00596387515808033, 0.0409662848299507, -0.0546100904677899, 
    -0.00685613139108132, 0.181778599236198, 0.12810939205382, 
    -0.00587047609381317, 0.0580056705275675, 0.355224927890395, 
    0.114144826656103, -0.00361373043675098, -0.128159807925178, 
    0.034789834249547, 0.546873047795173, 0.135617527579234, 
    0.00574384808746255, -0.283803749963932, -0.024296965231843, 
    0.704033382348255, 0.0972430010693002, -0.0727146118661538, 
    0.110771795469677, 0.590793784477322, -0.0991560696411042, 
    -0.0577799683654714, 0.102308719416198, -0.112270066121653, 
    -0.129644172165826, 0.0135748617479403, -0.138206126367885, 
    0.037092356031054, -0.119611953421083, -0.166538080673494, 
    -0.199263628961378, -0.143255776758918, 0.0428810872920279, 
    -0.169349876694133, 0.199150092774943, -0.164884648599053, 
    0.00751538215491883, -0.0760981319635776, -0.00223294828963708, 
    -0.232512425061669, -0.0194278402479725, 0.0366605126427663, 
    0.0709554062146461, 0.0822955131101775, 0.0898976447458862, 
    0.0631119584307251, 0.0567592493377953, 0.101834494817488, 
    0.0923213977244399, 0.0442122806640977, -0.0356137913727558, 
    0.100833477535149, 0.362247486903083, 0.193164998019932, 
    0.0593031275561675, 0.256901910916136, 0.177485395095155, 
    0.260936609009359, 0.498230985465744, 0.226652878996166, 
    0.0867466272947773, 0.0264464690550369, 0.0482646610263689, 
    -0.0574258803338305, -0.261948832800906, 0.797155945253726, 
    0.17481121747744, -0.202881796604666, 0.430444087077637, 
    0.529930004290157, -0.325859176676018, -0.0674763317493838, 
    -0.124271845558372, -0.0985780527730251, -0.0960332694436099, 
    -0.121738029697145, -0.0169533646003531, -0.134663102294738, 
    -0.136461382372177, -0.120987332980426, -0.153702353165289, 
    -0.0876590453638045, 0.0481355940016411, -0.0374259906511151, 
    0.15141456246854, -0.130679523307062, 0.0191640103366124, 
    -0.0768957791766617, 0.0111816906317329, -0.165164235635004, 
    -0.0185716371182944, 0.032334935219708, 0.0761797943063468, 
    0.0891919401778392, 0.078420729060205, 0.0620316796933713, 
    0.0924212485934415, 0.137501005770972, 0.0698948429001357, 
    0.136475035315689, 0.275286719437817, -0.137391358878346, 
    0.169992254952469, 0.561382378274615, -0.0191299125697243, 
    -0.0503503497456293, -0.181753736796797, 0.500269062376226, 
    0.247855468650903, -0.147301927194644, 0.506039915743943, 
    0.565213135092436, -0.127799567399495, 0.273145296238806, 
    0.600835031673498, 0.0950031537826815, -0.298958490973702, 
    0.403350084244001, 0.788777631184771, 0.182415945433916, 
    -0.0772078922495516, 0.0844579242139103, -0.152946529459552, 
    0.0602375377456455, -0.187755813953158, 0.00254722550954793, 
    -0.222117319837118, -0.0985782950071146, -0.0746024402529594, 
    -0.172558552664992, 0.0348904139117377, 0.0943623818754326, 
    0.0991569281182991, 0.173432481912146, 0.286427459684405, 
    0.28735384002061, 0.214469973937986, 0.167443468173616, 0.19062574930117, 
    0.270697563693477, 0.326490933331315, 0.255759367911724, 
    0.184061953492148, 0.294174870365589, 0.377485729441912, 
    0.213885242034228, 0.111620257444309, 0.408858146566498, 
    0.34968383623028, 0.110645365288282, 0.110665735238255, 
    0.501528432761013, 0.18926728099512, -0.15751464086457, 0.10698387035485, 
    0.62729421945497, 0.275416217996738, 0.0536838233437474, 
    0.113066004137817, 0.293514033663703, 0.696872920467002, 
    0.173171043879126, -0.213087212282603, 0.0137338163491245, 
    0.439716006084154, 0.0688494254755226, 0.29492716488671, 
    0.711245698981447, 0.248034798982618, -0.0286100972605837, 
    -0.139965705014075, -0.237529848152909, 0.0720214933224862, 
    -0.490385591042389, -0.143289140209246, -0.162979522004685, 
    -0.30641359255255, -0.129698254801239, -0.173287563263242, 
    -0.186508662402171, -0.0675303189360488, 0.110718227441827, 
    0.152816695912465, 0.155721321253858, 0.192158114125635, 
    0.189836093471155, 0.183975453492052, 0.208883100387299, 
    0.176000173520206, 0.135818482046914, 0.168208534435493, 
    0.174098675976369, 0.16307500935577, 0.236298221682848, 
    0.281786311854551, 0.180995354580668, 0.124790358913762, 
    0.346460574905575, 0.36305595912868, 0.14622149935473, 
    -0.127555754652314, 0.270903648081724, 0.464094146127257, 
    0.11716459521919, 0.0309658075723358, -0.215672375682776, 
    0.247910514590383, 0.446674146191603, 0.361369432308085, 
    0.101558420103536, -0.238398831462636, -0.025091729727751, 
    0.40254029116302, -0.0089496845087315, 0.624826309238342, 
    0.580656394642704, -0.074542696141675, 0.439103675524219, 
    0.696228639248237, -0.144839638165059, -0.104127641678474, 
    -0.126499871592633, -0.00613992642834432, -0.134462842682572, 
    -0.0258442215104311, -0.156154692840129, -0.089485708601971, 
    -0.1767500829578, -0.0636589343203747, -0.146432817776505, 
    -0.0517793824958485, -0.0210629167371394, 0.0239273541211715, 
    -0.00177711053957975, 0.0417615011074955, -0.0449697132159552, 
    -0.0528458829013944, 0.0488062893446728, 0.0238060876803889, 
    -0.082339111605037, 0.144750648305907, 0.194172843883326, 
    -0.168839331145055, 0.384350531919292, 0.29382893160556, 
    0.0377309396522253, 0.168140389629077, 0.367573561916692, 
    0.13814081449617, 0.209127717407907, 0.773740435840582, 
    0.101540748162955, -0.780833821289394, 0.264697050813355, 
    0.61749365885514, -0.348453005081544, -0.188191478609314, 
    -0.00290008445043545, 0.901775795798766, -0.107475712871251, 
    -0.0640208937831877, -0.00547634761084655, -0.0235301868754053, 
    0.201638697034005, 0.020053120676218, 0.018377429944581, 
    0.00902553943693529, -0.0392493800354452, -0.137761297965773, 
    0.0573138193092738, 0.253150243600971, 0.0976553788416375, 
    0.0672568821055223, 0.150406087426017, -0.027243114695351, 
    0.220756274090905, 0.0646100879079341, 0.0263838013734252, 
    -0.0532602593461691, 0.149885123587507, 0.123354068767219, 
    0.0396806302322125, 0.0101285033786389, 0.0170105070799232, 
    0.0518036245846242, 0.0713179608722924, 0.0949985686538719, 
    0.0224114555896566, 0.00103399093368813, 0.0105034808298426, 
    0.00409234092423945, -0.0579983974785185, 0.0250853184171607, 
    0.00591382114368021, 0.0272741654796925, -0.0379983640927213, 
    0.0222947491423789, -0.0327485405255984, 0.00748386094352182, 
    -0.0206494692276157,
  0.408506311055231, 0.302132970267527, 0.310543012801896, 
    0.0448048850920051, -0.0481700302224512, 0.0677073558608465, 
    0.18612569223522, 0.00329284881880977, 0.21014889251961, 
    -0.0258158871998853, -0.266273009170948, 0.0237299389812231, 
    -0.381924555366018, -0.162111944614326, -0.0736581513410241, 
    -0.363647744235819, 0.10738490613953, -0.0323382941221574, 
    0.0821841993858915, -0.241922942922809, -0.0629326764351038, 
    0.128494137315376, 0.22198140305395, 0.159766345191763, 
    0.136942742192942, 0.199206095207819, 0.2061293727213, 0.21525344587653, 
    0.276595987517301, 0.24076220814497, 0.108203812947476, 
    0.0670569665331021, 0.0901310456198295, 0.0594286351178673, 
    0.0794026160931665, 0.0999701042220296, 0.104140624032456, 
    0.0285346651932872, 0.0814418009744663, 0.0583460758821845, 
    0.0601495963293844, 0.0713433276616094, 0.0874414699479904, 
    0.081307919800208, 0.101227000549133, 0.108531539971836, 
    0.0679027933756308, 0.0821990601584422, 0.0635357642706033, 
    -0.0865014761744208, 0.167740394869096, 0.59411040107564, 
    0.157661384392976, -0.219960454474946, 0.0316659089724164, 
    0.562259689034859, 0.0659493116192306, -0.11201743668159, 
    0.167767703327502, 0.533819234901722, -0.0640452031058902, 
    0.0265847294612924, 0.162439640375263, -0.214478098448921, 
    0.152383524799263, 0.265985158281918, -0.0661250431963042, 
    -0.0401879743939882, 0.0151131329637602, -0.0786360978938194, 
    -0.11863111894144, -0.344898656859806, -0.081722183056697, 
    -0.0140690761867201, 0.0978364072183725, 0.00331126584532213, 
    0.163560559435513, -0.187841860223386, 0.0914079906889111, 
    -0.301532450102209, -0.0642456906617272, 0.0519317793409472, 
    0.0891351015244952, 0.0864911297453828, 0.132302049365418, 
    0.165972544797291, 0.169425987335973, 0.162077820824787, 
    0.120409770273229, -0.167782667479345, 0.48578055485625, 
    0.336929402526784, -0.0137178033164329, -0.0106636936370998, 
    0.577697892192837, 0.502448077564893, 0.204887453789401, 
    0.141630522427456, -0.295654956748933, 0.535082567649892, 
    0.328977907856632, 0.221262106908719, 0.653280029153689, 
    0.064190896995564, -0.385063086556813, -0.461234497404446, 
    0.954570144066049, 0.268842694840394, -0.147351702035173, 
    0.4565866646091, 0.410118731162668, 0.130153864226562, 0.055595653734211, 
    0.071875954376514, 0.118012110555338, 0.0964136008856119, 
    0.0840538232144136, 0.087108608556388, 0.0129866081573722, 
    0.0633889495532018, 0.358110824864115, 0.116560029093238, 
    -0.0550576464331743, -0.0570667366386127, 0.34252375816725, 
    0.290630810310272, 0.153883616995459, 0.0815548183642283, 
    -0.146093051916414, 0.137850321279982, 0.34411414615146, 
    0.0788901393853656, -0.0221372642180774, 0.523944071191057, 
    0.449666491471649, 0.234392259546001, 0.0696888977689118, 
    -0.21639711255796, -0.148537058996621, 0.623173332347622, 
    0.185362533035916, 0.0918063581086412, -0.160532994368519, 
    0.547558346958085, 0.255411756991428, 0.0827070257034548, 
    -0.103908274217898, 0.157658548833324, 0.278413832242398, 
    0.507857644494124, 0.310938576736309, -0.0828650837903207, 
    0.33262803027564, 0.372990453431728, 0.0793278241970457, 
    -0.0506247125920966, -0.0611082935896136, 0.546484337549332, 
    0.317221808786784, 0.0352182638281569, 0.426444800004333, 
    0.501912160808396, 0.207288880874855, -0.260680018456144, 
    0.432108766985174, 0.268455733066284, 0.014045677121072, 
    0.164933408429418, 0.509714379481559, 0.0368358417965816, 
    -0.0463422546450921, -0.0358876152203799, 0.000627298351866965, 
    -0.0344520132953128, -0.0043642809443047, -0.0347868013781997, 
    -0.00737767678534629, -0.00968354715968225, 0.0448765576789529, 
    -0.0951567322623442, 0.125955413278363, 0.189670813953135, 
    -0.0514601100398948, 0.16786399464859, 0.45938412389835, 
    0.0647530386313426, -0.0600750584959542, -0.121521338680074, 
    0.203950000879717, 0.401522047169135, 0.369679406373903, 
    0.156071461700236, -0.312607276879673, 0.155589054350096, 
    0.504249104090784, 0.220164360323014, 0.0855486072729553, 
    0.0584691252823523, 0.689405330911151, 0.116549712713766, 
    -1.0694097344513e-05, 0.149126130653281, -0.0299139449908076, 
    0.335367278558782, 0.112823415570238, 0.0416173046587446, 
    0.116864248443775, 0.254060041863957, 0.097983382559416, 
    -0.303181764767173, -0.269596399257195, -0.169786387584065, 
    -0.167657992020508, -0.264607110361143, -0.0907960203039098, 
    -0.282320150659769, -0.0728832765136344, -0.291097970583446, 
    -0.0827131431999107, -0.195715295174912, -0.0189685270131805, 
    -0.0701915658843662, 0.0253356558910522, -0.16207853215309, 
    -0.0529501944790937, -0.00827650548129144, 0.0193576742761752, 
    -0.038684584995149, 0.0220675843734175, -0.104701794251075, 
    -0.0285713629969507, 0.0498289333682336, 0.0753243840592976, 
    0.0751167277003353, 0.0856783073813634, 0.0891481294128508, 
    0.104767697985576, 0.127491974649697, 0.0818135940027223, 
    0.0093912084954025, 0.0631950992855501, 0.223523024539688, 
    0.212122345601037, 0.0671705253336199, 0.220407342437614, 
    0.441912958212034, 0.193993427806991, -0.0383777786881706, 
    0.250143246021859, 0.387601801896049, 0.200555828650431, 
    0.420100950024681, 0.485720398623882, -0.0647216734199153, 
    0.504452399428731, 0.403003431102826, 0.16415591355213, 
    0.550025714615381, 0.468366905841866, 0.140390164530754, 
    -0.049229762570939, -0.180851211889536, -0.0439798313924827, 
    0.101105910658721, -0.0759905991101319, 0.0238032210048967, 
    -0.114715795227033, 0.122105339813775, -0.043017061211067, 
    -0.0737162569687354, 0.0185154085311274, -0.272850301767938, 
    0.0739582218366453, -0.0956590856765815, 0.0666074800756319, 
    -0.205754810617017, 0.0350729105847822, -0.0747329809390995, 
    0.02883929151186, -0.283283624700853, -0.0395033935048635, 
    0.0654826567418438, 0.10560261182371, 0.195204042357163, 
    0.148972247167033, -0.0376102874939818, 0.126840083960995, 
    0.488223372863856, -0.0455749737285084, -0.201407592940135, 
    -0.150062833962216, 0.726375140201452, 0.0555853839559086, 
    -0.365677114715171, 0.119701847482152, 0.697805111408367, 
    -0.0368764644114382, -0.0914561380851069, -0.190277399228888, 
    0.527764116406711, 0.291048553074682, 0.0651288693892903, 
    -0.0958948061205847, -0.131988094787101, 0.215705970895689, 
    0.283929543306136, 0.395549226151843, 0.287765090016191, 
    -0.01666250750032, 0.279518575958146, 0.314982677551085, 
    0.00327797978397647, 7.79336919890794e-05, -0.101420976357471, 
    0.114573309066162, 0.0263889448760214, -0.00466976533973401, 
    0.125909176713184, 0.0352619789382519, -0.0687773316918072, 
    -0.119066564744497, -0.167462520584322, -0.0275279420559812, 
    -0.107300766429843, 0.000530087695360226, -0.178704905716251, 
    0.00711622670741143, -0.11722651483088, 0.0294026960692258, 
    -0.278473761927385, -0.021346035362524, 0.0651403322424666, 
    0.0534493069301738, 0.111805016727259, 0.183479240485449, 
    0.14582290518975, 0.118338167297105, 0.172643288949252, 
    0.160298955965436, 0.0842364689694893, 0.155196683838046, 
    0.270199808010541, 0.231672116842319, 0.119711980894095, 
    0.284196599018827, 0.43773691409763, 0.201499512160956, 
    0.029898167227317, 0.573138472090361, 0.260035243815427, 
    -0.0607505078256599, 0.0534065421899822, 0.524638377902284, 
    0.371604915846656, 0.198452824248683, 0.0790318049893513, 
    0.384078988936566, 0.13826410047464, -0.0868467180056596, 
    0.633932552309161,
  0.423078355003548, 0.436030767428657, 0.748297324585805, 0.133869433532655, 
    -0.20108384703752, -0.208102811023301, 0.939464595714809, 
    0.0303812631887367, -0.193292811656789, 0.416325365146033, 
    0.16166756676521, -0.0526519488656007, -0.0478255818817482, 
    0.0803345975587185, -0.159471017166537, 0.0920845265869349, 
    0.118733484909008, -0.0823321935620699, -0.13056083297363, 
    0.147814037906174, 0.0202529116091937, 0.101822790640302, 
    -0.0291089561071245, 0.11579942055962, -0.185770991784431, 
    0.0348489699667553, -0.343774030898349, -0.145557278347091, 
    -0.0379893256891489, -0.210170623234351, -0.0100874038663862, 
    0.0422109964113805, 0.114549007240206, 0.159392561185277, 
    0.164371338434849, 0.1699146475469, 0.185974163084952, 0.179585516420154, 
    0.146168654411897, 0.144303854796425, 0.237779422022174, 
    0.243486569136459, 0.195167623125077, 0.218582415901613, 
    0.308325210612293, 0.258838151885439, 0.138082924488475, 
    0.147146965995647, 0.356567732405825, 0.323545739884965, 
    0.142454196855812, -0.0833205098735507, 0.152701243736949, 
    0.460423135372739, 0.234852607516605, 0.110974331302274, 
    -0.157317905504937, 0.402109645174287, 0.358729814959561, 
    0.15998224968134, 0.0254993181191923, 0.326091941011305, 
    0.201527840204179, 0.0457795164767197, 0.150361590126282, 
    -0.388591151225676, 0.596433332367742, 0.516950305363581, 
    -0.347239927970292, -0.165224751713937, -0.310073531207518, 
    0.00729855731055967, -0.311513947797699, -0.0998923739106146, 
    -0.235892859411255, -0.204726814879748, -0.0156909857710134, 
    -0.238805776790749, 0.0789358035549262, -0.196205573737737, 
    0.105115366170644, -0.0210719345947131, 0.0662158754093761, 
    0.00672273750899367, 0.0738393239750206, -0.0378442882129416, 
    0.0515488607607079, 0.0160640330002446, 0.0781776412241608, 
    -0.0223638792503214, 0.0665391868569758, 0.0340295225252062, 
    0.0357807982242045, 0.0369397205536463, 0.0404006132830833, 
    0.042977420629247, 0.0480936349527834, 0.0521601888236241, 
    0.0577289836469244, -0.0142291440184967, 0.145964446382249, 
    0.13841451756974, 0.0496975628015572, 0.263456443832023, 
    0.244625359752551, 0.0486191325406035, 0.182430207371159, 
    0.358144110981815, 0.223480200588182, 0.159048585037895, 
    0.080624487525387, -0.276117903366124, 0.02954986403445, 
    0.659153713199652, 0.131126106560308, 0.0250387186637439, 
    -0.300278687942924, 0.173467264903917, 0.589009121468598, 
    0.254613240302899, -0.0117663726463883, 0.288648976852983, 
    0.151641455545043, 0.117060160121238, -0.378066055240268, 
    0.189609561687693, 0.185005754838888, -0.0777062914328382, 
    -0.10852604617944, 0.272772359734959, -0.100084423740194, 
    0.154049498455541, -0.25403703439705, 0.0757295308685814, 
    -0.162295430679932, 0.0400038457884402, -0.385995194991967, 
    -0.0331122067429447, -0.39907760819204, -0.242390381972264, 
    -0.0468016984829402, 0.0582599134227198, 0.00671067372403675, 
    0.0334420064983431, 0.0294945504289489, 0.0396398703500325, 
    0.00720862549034937, 0.0411673330671282, 0.0603557853846768, 
    -0.0898952007945898, 0.332161953245045, 0.26792080848995, 
    -0.0775389394200491, 0.202618936516376, 0.455404798908597, 
    0.140682020802055, -0.113153567703986, 0.360183825614639, 
    0.553582634497453, 0.431841418613854, 0.251821684596298, 
    -0.236182725734306, 0.252473580870715, 0.37477804113672, 
    0.11220167920322, 0.881264419296895, 0.467789270645312, 
    -0.101155150948177, 0.474667225722616, 0.491974933816134, 
    -0.254715020469197, -0.273717071333194, 0.0307644670505082, 
    0.288857363631576, 0.0927354017267083, 0.0378028725858516, 
    0.0480669959165481, -0.122218607334696, 0.274124766155971, 
    0.169782838435618, -0.0809141909200036, 0.137638507658979, 
    0.389446420892949, 0.24427938817437, 0.116911617856332, 
    -0.128271845543022, 0.179449874859449, 0.268759677553507, 
    0.114910850092519, 0.0357275828029373, 0.0300857428611709, 
    0.205812888651423, 0.158451468778426, 0.0488226202997043, 
    0.0143877675942074, 0.226699745647931, 0.157465658781228, 
    0.117036065336084, 0.11003124626881, -0.00667138769250112, 
    -0.0787129820192426, -0.170843199542566, 0.0577422210409179, 
    -0.105178487383391, 0.0543517676050045, -0.161507142652519, 
    0.0594465968833723, -0.124315512307472, 0.0519139929323859, 
    -0.207411965633335, -0.000325692112563947, 0.0455084303624954, 
    0.0682451373772161, 0.116840041116953, 0.138901729127294, 
    0.124528531938142, 0.143779990655624, 0.156525965641325, 
    0.0882946334825349, -0.0394751645834261, 0.357962373475207, 
    0.276369370775818, 0.0763695135259675, -0.101838664536995, 
    0.428700249209591, 0.360757208809712, 0.113706163189471, 
    0.0698767503199603, 0.469427992892475, 0.248850465155689, 
    0.0461252624308936, 0.786746402815624, 0.252472112374805, 
    -0.0483008620031143, 0.113408468938713, 0.635609061346257, 
    0.0359249070253925, -0.323402028206279, 0.30099741448888, 
    0.354237871556213, -0.188957756738537, 0.00343092231314512, 
    -0.146728898810651, -0.0405727319211897, -0.10967743980672, 
    -0.156911188256397, -0.0780074123181851, -0.107562953748012, 
    -0.22927342113429, -0.0893711764302652, -0.0841247364309379, 
    -0.109151529192029, 0.0537112389816921, -0.00856233692832382, 
    0.118472461412893, -0.0678438047900741, 0.0378189117249522, 
    -0.0340604105565531, 0.0529182018658684, -0.161969226981979, 
    0.000273616448288577, 0.0649047432254137, -0.000167587794095023, 
    0.105290033737937, 0.142175836282529, 0.129147505997771, 
    0.155418599430181, -0.181436182502307, 0.31039307885325, 
    0.18023558917582, -0.0626286574162822, -0.0128463898905797, 
    0.598748705576533, 0.415986193886578, 0.25395687049624, 
    0.153345868258982, 0.185516936491817, 0.470030945538984, 
    -0.367253857715427, 0.168164103993548, 0.912888347254141, 
    0.382092458889522, -0.00188467047981708, -0.271282660087781, 
    -0.462266951340615, 0.388003230797205, 0.701018142678774, 
    -0.0296320195534088, -0.030480678234214, 0.123132330630454, 
    -0.607356170210168, -0.039289524044434, -0.487441408639064, 
    -0.319385774727531, -0.0744476728618097, -0.390544763508398, 
    0.139781435546192, -0.333603887869529, 0.144535071605666, 
    -0.40233449654134, -0.00112047657863985, 0.0471456286073904, 
    0.0761809561233903, 0.0674974564047152, 0.0921361340222512, 
    0.0705596203698183, 0.00127199577099338, 0.114623303776726, 
    0.156640020234602, 0.0853114629674685, -0.0330833212525617, 
    0.224794882170939, -0.0660025127115857, 0.322882524885577, 
    0.851054958918439, 0.0416587622740007, -0.039089397421881, 
    -0.068720210215738, 0.64421644772081, 0.140917824253917, 
    0.018269250297901, 0.0766957692561193, -0.209333862310188, 
    0.265657995456834, 0.205830814203471, 0.0571320347230479, 
    0.355764373785754, 0.191029063603159, 0.0194347626820382, 
    0.0165238676393265, 0.0326682670217744, -0.210170722715572, 
    0.153501898099638, -0.158801012623789, 0.0600776238341714, 
    -0.25956610991488, 0.0186331185206278, -0.146847856548945, 
    0.043541286561736, -0.316832907511915, -0.0319872058331928, 
    0.0654642616723099, 0.0846216014510157, 0.148591719909844, 
    0.180048465285495, 0.127006334935968, 0.11837492785626, 
    0.214277885186593, 0.160899109573677, 0.0334139072228573, 
    0.0600098448116851, 0.331638822745394, 0.291382273823957, 
    0.157816867836943, 0.160949123268331, 0.221146894512483, 
    0.460010301477213, 0.328685893288046, 0.0352055464904761, 
    0.341171647551691,
  -0.106946135985832, 0.0394119013472882, -0.216834220376025, 
    -0.0691291667160365, -0.0687666403256007, -0.0935444500406404, 
    -0.116214129991862, 0.0751434391894395, 0.0201525891729284, 
    -0.0841601935594026, -0.265336013351207, 0.246319153804035, 
    0.277665016318879, 0.115566152806517, 0.498166089165132, 
    0.372677318624174, -0.0907083420827294, 0.345686670136204, 
    0.424097079671679, 0.0537428974186926, 0.160739153830317, 
    0.719606581242364, 0.0437487434906471, -0.112752931200312, 
    0.107511755713912, 0.520708607918348, 0.0356376348166695, 
    0.465554286446308, 0.641326133197202, 0.0268255791694533, 
    -0.0752817742869529, -0.0591984094797524, -0.0109356680217497, 
    -0.0716847254137505, -0.0179095026313586, -0.0719071514096463, 
    -0.0275171096980121, -0.0508719621398689, 0.021548602840928, 
    -0.0873207895126807, 0.272046519738194, 0.0991403420251892, 
    -0.0655629765432738, 0.0219142457685908, 0.406240908321296, 
    0.265234808364646, 0.105870245902893, 0.0819979114761373, 
    0.00255204246949259, 0.584753655780958, 0.286655023193156, 
    -0.0343224093171253, -0.0262082164794814, -0.265532565531314, 
    0.468710936426623, 0.300049442136686, 0.114023808056747, 
    0.425073206462351, 0.406641352043639, -0.260320954236741, 
    -0.223789121936946, -0.119241520976876, -0.13119445302465, 
    -0.245553593417927, 0.133816887349117, -0.155781519731869, 
    0.0358384567274563, -0.0755792292715961, 0.0429391567215561, 
    -0.222706684235622, 0.00726487094811881, 0.0984846425830976, 
    0.119908997391837, 0.199468005770748, 0.272136103765591, 
    0.219878689040193, 0.155862855665331, 0.180526512615878, 
    0.233247241471429, 0.226853485444313, 0.211442663613094, 
    0.194278373646429, 0.183863876800438, 0.209322324126024, 
    0.227272894432908, 0.184572400967829, 0.162275458032942, 
    0.242890849607826, 0.249935264586545, 0.168136612623761, 
    0.165205884181481, 0.215298174377192, 0.165501826924471, 
    0.243101126530742, 0.358613182905936, 0.175447528032048, 
    0.0382385120177684, 0.493461021621704, 0.337276121603395, 
    0.0534138616778893, 0.0950478105595265, -0.310360060193884, 
    0.336549329479689, 0.308742567771431, 0.145705150550756, 
    0.645476864260323, 0.349188406299034, 0.094022415898622, 
    0.581761962851247, 0.163289324652325, -0.259763374910822, 
    -0.0914231958246263, -0.0853169333110462, -0.147652614984366, 
    -0.0397282846747951, -0.236200010092433, -0.0897281488352773, 
    -0.195034600856862, -0.0290706508532687, -0.172060047449705, 
    0.0424256656365658, -0.216004741520965, -0.040765774038638, 
    -0.0343410945696894, 0.0525254601709934, -0.132057286757268, 
    0.0372526101185368, -0.0341088447896841, 0.0376701775910036, 
    -0.23822631365593, -0.0541701178388643, 0.0960878635454916, 
    0.0565685637753373, -0.0696356851496182, 0.0638708101699545, 
    0.218614203114003, 0.094199364538155, -0.000428241230985088, 
    0.120846483312515, 0.261140579388653, 0.278690962449931, 
    -0.281133659314855, 0.568589885664282, 0.665423969342053, 
    0.141839274725657, -0.0698337545101861, 0.00445025150241056, 
    -0.11413973969748, 0.371000525041374, 0.892288705726045, 
    0.324278026945005, -0.0518903432631756, 0.294302800493468, 
    0.169518490747115, 0.779396715948146, 0.640189865293336, 
    -0.0269536185819675, 0.132156163970661, -0.192746938210317, 
    0.628333594258863, -0.0539687144112236, -0.116339955248224, 
    -0.152526771284336, -0.167194250116353, 0.0753831890505888, 
    0.0299159632895686, -0.066823703497812, -0.132254886036868, 
    -0.0892142193145627, 0.0427170248650949, 0.0897369562349571, 
    0.0581346882292647, -0.00841170064814743, 0.0954684931091017, 
    0.0903231922060286, 0.14252233116939, 0.255004801838393, 
    0.150248844231067, 0.0134951658978546, -0.186275063267887, 
    -0.0128257174342617, -0.0121986653905043, 0.927169937020694, 
    0.0934633799153895, -0.108253400223773, -0.451248895954933, 
    0.535090040969234, 0.691352520108179, 0.279005105216925, 
    0.279241008983357, 0.702730979169253, 0.020735011554657, 
    -0.151990185470324, 0.227204506730365, -0.119609522241573, 
    0.304538766426538, 0.222361924436583, 0.751772014844064, 
    0.35945307014583, -0.0799065516642784, -0.0891999192693529, 
    -0.0719648397081282, -0.0891752382211686, -0.0705568528788407, 
    -0.0854791676228669, -0.0199503021898671, -0.110560556638621, 
    0.0190300247314981, -0.0726792802268219, -0.0238777185716861, 
    -0.0484719993796492, -0.164572390304183, 0.308537050512769, 
    0.410127908553021, 0.111591644757282, 0.0117237829340814, 
    -0.267482177773613, 0.0406346719228925, 0.544589942711474, 
    0.262746560922729, 0.025122367245546, -0.00924711633437451, 
    0.391700922586234, 0.164282373714181, -0.00561201667351832, 
    -0.0122323674612113, 0.269975818784676, 0.285359274550289, 
    0.164155346253331, 0.0505684630914134, -0.0471221283413647, 
    -0.0984040943621064, 0.107686203005187, -0.120871653792026, 
    0.0108497615638473, -0.174827234227365, -0.0519790213309884, 
    -0.0983334561494354, -0.0585034284480917, -0.126222272419067, 
    -0.106869870939955, 0.125810046226794, 0.150705836521649, 
    0.0611270234185026, 0.0189500081860992, -0.0129765461867, 
    0.330605558665811, 0.245646769026996, 0.0239126089376683, 
    0.100873862064534, -0.324734938880798, -0.0580268641381198, 
    0.515961902920238, 0.351106029097685, 0.280773599800328, 
    0.53917827639182, 0.240043169727677, -0.165835457560644, 
    0.981242818939601, 0.407895068910871, 0.0828541570694378, 
    -0.244008957761685, 0.233184726645328, 0.775986189715019, 
    0.398985866404144, -0.0761325142711127, 0.64618861421378, 
    0.738772324606516, 0.363681817551783, 0.200266067567602, 
    0.124107056376809, -0.251066416882821, 0.420808637851238, 
    0.321865722973428, 0.0298893079819127, 0.174220525969317, 
    0.279082095709794, -0.367075197897427, 0.198449237412046, 
    0.186311097720888, 0.00807427558679983, -0.04835295050059, 
    -0.225222380359248, -0.177446848358657, -0.144507709831599, 
    0.0840304065840908, -0.189921277236217, -0.135733668299741, 
    -0.030262230118607, 0.0704698231410727, -0.096577160991563, 
    0.00466020961340967, -0.115557148266058, -0.0466169807092072, 
    -0.0602031217883593, -0.0844272019058961, -0.0151917975334122, 
    -0.0890148390786674, -0.0421215945292723, -0.0116258953520614, 
    0.00295119020154935, 0.0537663939327751, 0.299190535247421, 
    0.122625393032447, -0.0513778124969203, 0.395808157476522, 
    0.396621766415033, 0.192781543081699, 0.0804892615393506, 
    -0.195120462667813, 0.00711550161905018, 0.432883612141531, 
    0.132753934404377, -0.02640889276407, 0.111366753484744, 
    0.24964306418217, 0.0744545608050796, 0.342001320898682, 
    0.390521346406133, 0.0401844956509648, -0.069908378354193, 
    -0.0165514365685272, -0.0639116479328676, -0.0448208966734717, 
    0.00523755162854236, -0.0445975731837568, 0.0177799353904449, 
    -0.0377319689502676, 0.00778461691488643, -0.0661413143762802, 
    0.00916518496065427, 0.0709435426768347, 0.114508498246642, 
    0.0931333063704251, 0.0550702336686169, 0.063141827605812, 
    0.19210176653752, 0.145329181204022, 0.134575142572223, 
    -0.247044946493153, 0.437701227415046, 0.323107988334014, 
    -0.0719838623736595, 0.859326105313762, 0.539886405053543, 
    0.0985908490728404, 0.299807032848864, 0.0325970526487744, 
    0.996373997971972, 0.04646022330912, 0.0141994810935392, 
    -0.226329785067447, 0.0713843451243441, 0.19932742758584, 
    0.0111636975005977, 0.00507022664501046, -0.109415345416512, 
    0.177224434315393, 0.0829147311825371, -0.00811236666511642,
  -0.186222260366433, 0.110198360280233, 0.662584677297313, 
    0.253393942082546, -0.0343651755084905, 0.288913321347472, 
    0.312682790782902, -0.259386249805496, 0.768152711575021, 
    0.509629516007764, 0.0505841175767893, 0.0293629762575097, 
    -0.0206539813256876, 0.0355262469072867, -0.0387633436238082, 
    0.0120582628740362, -0.023855833774985, -0.00938939363204219, 
    0.0253265577522623, -0.0429282231289122, 0.0403417938102592, 
    0.0833891914606232, 0.142357151491647, 0.16638533677103, 
    0.150868538302923, 0.120941065488297, 0.172762789047388, 
    0.269699912105337, 0.159093424134898, 0.0196142413966729, 
    -0.0290994552142413, 0.392277776598758, 0.32863456886869, 
    0.112217559742453, 0.277391992565141, 0.390032425162375, 
    0.0769794715996949, 0.182354263546966, 0.377781594912429, 
    0.455670796814862, 0.780109837541487, 0.263954392040001, 
    -0.0781855604858921, -0.411740075012505, 0.20265246118819, 
    0.888280487947573, 0.127664290064378, -0.125872223953859, 
    -0.15403300900297, 0.5898619531381, 0.308287409376375, 0.262410322318142, 
    0.24899344326924, -0.029369024419153, -0.071647271690106, 
    -0.20529103689641, 0.37912312259332, 0.100574015641127, 
    -0.116094445408537, 0.167572472659518, 0.290956452060255, 
    0.088045343834508, -0.000670443758120975, 0.259581018637286, 
    0.193163618567821, 0.0790441453054074, 0.0465944664590385, 
    0.0570915105789456, -0.174192416847, 0.0517851588170728, 
    0.295491155164398, 0.416011295780671, 0.300804216666376, 
    -0.210463897455677, 0.294551956212225, 0.491526423689158, 
    0.260172474533618, 0.122489230034206, -0.0362054326645553, 
    0.117389430090166, 0.556594638047648, 0.0822777698259506, 
    -0.0261759148569078, 0.0720902829104705, -0.0688583336448158, 
    0.189035846383585, 0.0737520756735901, -0.0458534672501031, 
    -0.094577995758663, -0.228434954145417, -0.0136406441054486, 
    -0.191067411788067, 0.128190590284776, -0.199305810357845, 
    0.0503912193963201, -0.0781301471004602, 0.0617049055633107, 
    -0.255739887194334, 0.048430468905201, -0.121689092776303, 
    0.119805052875387, -0.0374943161067873, -0.00213518654929946, 
    0.0470341765211189, 0.0680711797125016, 0.101674768579472, 
    0.0184810233261203, 0.040439864812979, -0.025859880421275, 
    -0.00589033639501551, 0.0464205999367597, 0.048170281872063, 
    0.0570001034049229, 0.0413686313508759, 0.0562595943933377, 
    0.0526870588743615, 0.00566143545021931, 0.115411245029831, 
    0.107436552275493, -0.106966717619476, 0.152644785691753, 
    0.29125303053781, 0.0780102933187974, 0.120153005087136, 
    0.237292181202687, 0.0616430349978789, 0.144334540498157, 
    0.399378741410972, 0.693507894450841, 0.385267319963669, 
    0.0610238531687921, -0.229502661610427, 0.516283863466637, 
    0.549820214809936, 0.220561788326974, 0.0633932680555493, 
    -0.468354093176681, -0.313199840772506, 0.569226052442718, 
    0.336437553790713, 0.0218373430688457, -0.00271097659257985, 
    -0.243355157868506, -0.203841488336771, -0.243174217469385, 
    -0.1784719244155, -0.198965166793714, -0.205817112748753, 
    -0.0174631950964462, -0.26607449003779, 0.122631836385469, 
    0.0152047263323825, 0.0989263786377606, 0.0174821679640478, 
    0.0923106964017514, 0.0252236008399265, 0.0799227324132378, 
    0.103420298450993, 0.0888144949674048, -0.0504995851283018, 
    0.0272093850274881, -0.0581737397825572, -0.00193775260077596, 
    -0.0347720243816942, 0.00614962433348289, -0.0475061905442037, 
    0.0178219961122862, -0.0314868024121076, 0.0469633742296328, 
    -0.0690921310560024, 0.0515871543623702, 0.0878581360885918, 
    0.0948158431961638, 0.106449842474094, 0.109359216030612, 
    0.0980650683106808, 0.0811388856048154, 0.0728735088072837, 
    0.135304276791082, 0.116248629048208, 0.0155070481533662, 
    0.00879845128778206, 0.0520754537747611, 0.0136395617063906, 
    0.0344357708025079, 0.0195719784587782, 0.0382342002177605, 
    0.0598489087122467, 0.0863833033439535, -0.0503077299120409, 
    0.00403126369329035, 0.168951686823029, 0.255424290466238, 
    0.149718331002811, 0.0969835896650518, 0.205660672572935, 
    -0.097331480414541, 0.546158610992305, 0.167158811333394, 
    -0.24081448524082, 0.374418946735251, -0.0386213218033562, 
    0.857692974265333, 0.190521213342809, 0.0667546986762287, 
    -0.140434608325008, -0.250036870424032, 1.00848372273031, 
    0.758069886563908, 0.278239531238915, 0.118725131508043, 
    0.212416113354822, 0.130001676328587, -0.371773294380101, 
    0.144628032039584, 0.542708057684652, 0.0755483044457252, 
    -0.227082796453172, 0.0793874394119809, 0.654628276349421, 
    -0.00158973824746384, -0.129708694346867, 0.0931669071080955, 
    0.294768021650637, 0.0336360515062214, -0.152054372422715, 
    0.0923311769515187, 0.431576604148331, -0.0201610223237707, 
    0.111727077825594, -0.296223695998684, 0.224682031223282, 
    0.462461185185197, 0.0929251053900409, -0.0369155059356777, 
    -0.210549768612142, -0.0564899303851914, 0.706710975674672, 
    0.18300822395182, -0.0902098171849488, 0.0240101529930496, 
    0.373851994075897, 0.349780570468211, 0.377436538028587, 
    0.281815934469524, -0.159183749548181, 0.72171785389059, 
    0.404925742875619, -0.0337835439994083, 0.0478278195460885, 
    -0.34358461066361, 0.392765472995997, 0.402853231586024, 
    0.220222992661908, -0.00382512365270637, 0.514047079905981, 
    0.228208244591634, 0.116677528434669, -0.0992371943148606, 
    0.358740244292991, 0.236605254403269, 0.101412941584536, 
    0.0956886849552683, 0.119574833586509, 0.0477222947513621, 
    0.341140124378099, 0.045544934165034, -0.020590893025743, 
    0.0101795840228367, 0.21892369341794, 0.0850834439472874, 
    0.045679282376518, 0.0532841832939482, 0.0805112316866898, 
    0.109286403205831, 0.079756812208534, 0.0305930512984664, 
    0.166417142231366, 0.0403504024390999, -0.00078915332677458, 
    0.043202210941576, 0.301712479348632, 0.00626242978526366, 
    -0.0933984949824856, 0.559376413722274, 0.561313078557565, 
    0.0817762531655161, -0.189948658586628, -0.104722282627191, 
    0.348743687362316, 0.328349112721893, 0.222186212123959, 
    0.0655771977487426, -0.0595553853720113, 0.0686542419225722, 
    -0.00122219895777827, 0.246504384296369, 0.400626646816544, 
    0.131896884144801, 0.0064763274665172, -0.0490374132744604, 
    -0.129732468523203, 0.0538634146987516, -0.103849828297023, 
    0.0431877716632226, -0.152572451521327, 0.0230431095892151, 
    -0.174614787108824, -0.0326159495641144, -0.0996678252121308, 
    -0.00640207547343841, 0.0623635662287888, -0.014072796861404, 
    0.164887862693114, 0.0882532985539266, 0.0781998531212783, 
    0.180068906362495, -0.220168185893034, 0.247884592809496, 
    0.594165405148234, -0.0956581979055082, 0.19682622423843, 
    0.589652526859617, 0.193612112116527, 0.875443316991888, 
    0.825045653435021, 0.187201544027519, 1.00653688479834, 
    0.0255288232559066, -0.499804765950817, -0.17164755159718, 
    -0.154768318317193, -0.0534914651337483, -0.173894588926919, 
    -0.0390996721832463, -0.17289722987973, -0.117963633842842, 
    -0.00362750422614133, -0.1291219578487, -0.0496405724497165, 
    0.0570372494071, 0.10331659389148, -0.00735421448874425, 
    0.0167808237306233, -0.164757984679742, -0.056547388696718, 
    0.0583731529227148, -0.039263570295667, 0.085025584163457, 
    -0.119461647530794, 0.0292940627499676, -0.0132163751155763, 
    0.0691464381852309, 0.212550178053684, 0.101534889978567, 
    -0.0773332996825307, 0.122079337761374, 0.278191438460994, 
    0.0213130337057194, -0.0863022892394361,
  -0.0359758352110644, 0.0871807031373134, 0.0934735030002263, 
    0.131854883926636, 0.0155796168548586, 0.0891886446149612, 
    -0.0665162064381436, 0.0244720851879624, -0.0248475156614932, 
    -0.0294060939079149, 0.0244561954145753, 0.0691376465571159, 
    0.0678969860491893, 0.0723620747568972, 0.0782307127643926, 
    0.0641903719337731, 0.0788680729947564, 0.105841349634274, 
    0.051800148024544, 0.00676926290402614, 0.12254921563491, 
    -0.170508044419412, 0.266958817643324, 0.469555344888176, 
    0.149407151058883, 0.0016374682477851, 0.012563085677149, 
    -0.364561497464497, 0.438034678533413, 0.322069522622087, 
    0.318960860342141, 0.405636273973612, -0.0393181831271686, 
    0.749833331866858, 0.660257098767623, 0.286225203349755, 
    0.144713213046385, 0.370545904496746, 0.762163152483065, 
    0.108098631376241, -0.0708117703545175, -0.1174723389981, 
    0.0605693834147715, -0.00879259732619162, 0.0263474196582136, 
    -0.106798440857798, -0.0132455718482094, 0.0140431460153483, 
    0.0318065359725307, -0.0946632410468677, -0.155765113772795, 
    0.264545624326505, 0.319454977216842, 0.0903610873047683, 
    -0.183734379187073, -0.0333930618497023, 0.457769826472447, 
    0.315164961571406, 0.143061657121093, 0.0581480683717818, 
    0.0350943293730779, 0.112327411011205, 0.216992218629626, 
    0.40303895569703, 0.567923136298509, 0.466541203354459, 
    0.236399675195296, 0.0568504290666094, 0.35258582268851, 
    0.590961830102958, 0.263588454713836, 0.0516744502364547, 
    0.386005275878178, 0.369991402779408, 0.0351790178397587, 
    0.161135732787118, 0.561424965099123, 0.258159890626184, 
    0.0447604556576449, 0.402153769465253, 0.456942817628247, 
    -0.14122118911082, -0.349887723292787, 0.293347302512635, 
    0.200804677609498, -0.338152640655147, -0.342356554444171, 
    0.152269502419614, 0.444249860908819, -0.282602405733516, 
    -0.120978836463864, -0.145977328061636, -0.0631355520025356, 
    -0.189825109385384, -0.011926365242272, -0.281064360410322, 
    -0.0444623680307841, -0.216447971994737, 0.0280763179536119, 
    -0.134976872418491, 0.0996618662776414, -0.10069299814852, 
    0.0238527597848297, -0.0166127992662816, 0.0493107418368851, 
    -0.0774380763196529, 0.0482218656379739, -0.0877898884312915, 
    0.0258894362055659, -0.163291147014639, -0.0225623174896769, 
    0.0498598446855472, 0.0762240561390156, 0.127774588348279, 
    0.184471824810172, 0.131843777823255, 0.0620483683365573, 
    0.0341951413794587, 0.10275427910025, 0.370141165872205, 
    0.368378039931501, 0.168337465604328, -0.31297382910811, 
    0.388978796797663, 0.45614849399726, 0.0438838883101735, 
    -0.00119210183719398, -0.29497898139665, 0.451897392409777, 
    0.322477542387638, 0.166870430517024, 0.389039319574953, 
    0.231213386212233, -0.391604432051915, 0.256450880439552, 
    0.430903370868236, -0.0133014765117126, 0.127220504915464, 
    -0.148191603000256, 0.435758787606688, 0.0893089466963217, 
    0.0109608069850709, -0.111329566372523, 0.0936780462785986, 
    -0.0912012385581812, -0.00903461053455086, -0.150544792433037, 
    0.120408172450767, -0.056825276617463, 0.0718635419900916, 
    -0.114999626276288, 0.113990897778205, -0.207309601831164, 
    0.00882118254574671, -0.0883024178324197, 0.0372315224873137, 
    -0.225873324397236, -0.0217408042874208, -0.293272373453723, 
    -0.193439363600991, 0.0353630561755303, 0.0125950356627817, 
    0.0783927958238041, 0.232170559168467, 0.231203159245913, 
    0.087375827478185, -0.130323618879978, 0.035430666161879, 
    0.288030740741462, 0.368692309708299, 0.33554484561915, 
    -0.137332589838055, 0.649651854134068, 0.592609055276903, 
    0.0241846593029213, -0.0741801274185462, -0.339138003607355, 
    0.777867047258382, 0.203054055876794, -0.067432334221168, 
    -0.0782041732638874, 0.337764594482855, 0.475470787340012, 
    0.392467387741505, 0.247904946957309, 0.657867937142706, 
    0.587190720935786, -0.268837900786315, 0.576986324900585, 
    0.619456296348269, -0.203714024982833, 0.019888155873546, 
    -0.237307720698247, 0.242400122658917, 0.361404866419792, 
    0.0651006606032115, -0.481300642922539, 0.166176411136812, 
    0.248088320128135, -0.449969475439967, -0.198700495945719, 
    -0.038540542776768, -0.142234419702542, -0.112081612167549, 
    -0.105910744062173, -0.121397843207168, -0.067866071371134, 
    -0.124047656672037, 0.00675249841304065, -0.1635214111048, 
    0.0347457040936829, 0.128320863131907, 0.030177414882722, 
    0.125042613487291, 0.355307392762673, 0.151155886229761, 
    -0.0292836863869729, 0.0147572138576883, 0.444016584103152, 
    0.194953341018248, 0.107461505901722, -0.211169870081455, 
    0.00500301236271666, 0.71356113383872, 0.208280840647207, 
    -0.00366141734667971, -0.0749494715769539, -0.119309598649466, 
    0.756428717566825, 0.358523523730564, -0.0347946164011283, 
    0.388857582037987, 0.412501530343564, 0.0986723929754551, 
    0.109955203994435, 0.457981692938654, -0.1085095643891, 
    0.165900259832782, 0.938705654804765, 0.140519452186601, 
    -0.0917036514189255, -0.226989510815724, 0.0180452985478918, 
    0.0975763677224485, -0.0131512713852276, -0.107849921453734, 
    0.0401642551201397, 0.0704022512325992, -0.0358377079755552, 
    0.148463812154093, 0.0133322836000847, -0.083875350530689, 
    -0.0472808115946974, -0.0796462641694215, -0.0397918178948274, 
    -0.0145305923296716, -0.0423984516096939, -0.0101247361022986, 
    -0.0670724671909682, -0.031552411911544, -0.0155034602241955, 
    0.0454603168046115, 0.00629627517054655, 0.0350211236474706, 
    -0.00712412856583955, 0.0194002523566642, -0.0369485419045243, 
    -0.00980098954359807, 0.0319211901021273, -0.0100028767187551, 
    -0.0428781822736645, 0.211392045811976, 0.186199440967031, 
    0.0349810448341577, 0.0966557263099592, 0.202213425541468, 
    0.379503715948968, 0.317524795646572, -0.0417134452518427, 
    -0.07522581964165, -0.36597541072933, 0.131191899807873, 
    0.619013559426241, 0.157433810692894, -0.18707844674278, 
    0.100574095798616, 0.469121850366666, 0.0566417173998796, 
    0.439917014335458, 0.752507209050658, 0.0689875504952784, 
    0.0285449244462437, 0.0747959930415283, -0.0647024370916624, 
    -0.0721185059382485, 0.0310104469406427, -0.0133667845220755, 
    0.0468955976805927, -0.328437372391207, -0.00535248730034662, 
    -0.274097575667155, -0.0734477227940132, -0.20631569586086, 
    -0.170496313287273, -0.0377447991033122, -0.178567322585979, 
    0.0647905830643433, -0.147432411931329, 0.0918406696953125, 
    -0.10136657995727, 0.0994099714142832, -0.0311044309637873, 
    0.0165128416750787, -0.0138073032442856, 0.0186996118421092, 
    -0.0162701506954176, 0.0239093602921298, -0.0277172470763846, 
    0.0385332396752215, -0.0719169976656254, 0.0490381579171309, 
    0.09128469174029, 0.0320037942639679, 0.0767696676745911, 
    0.210268549030914, 0.146282755933227, 0.0806544025531167, 
    0.110092119195771, 0.208020321464239, -0.29838609065919, 
    0.441251045792301, 0.395620306092389, 0.232151612430168, 
    0.183253200245244, -0.296747644235586, 0.515118306242219, 
    0.495793284994476, 0.244126206461396, -0.12329003066321, 
    0.471720255896166, 0.300299026001094, 0.038925744194936, 
    -0.0221852448253414, -0.123533204179406, -0.124479622415465, 
    0.36064660303405, 0.140034666018318, 0.0657979707352882, 
    -0.0354510790031426, -0.331711031867305, -0.431920800316005, 
    -0.164101733485022, -0.192653663102037, -0.345638306148641, 
    -0.10783655670324, -0.337911169333395, -0.232302239727379, 
    -0.185667980227969, -0.247626019078751, -0.225180308394093,
  0.388806509356791, 0.0486632600824683, -0.476062405494717, 
    0.546006547102266, 0.608835665420812, 0.342251622733569, 
    0.343822323833899, -0.335456395160379, 0.508621395157009, 
    0.197138600103341, -0.114982967189068, -0.0435703047625847, 
    -0.129797369578395, 0.189628934928773, 0.052253390548675, 
    -0.0583163438274342, 0.151626351044094, 0.0983921723646418, 
    -0.245305667651243, -0.0635112835796714, -0.29540931719673, 
    -0.174368735315915, -0.102347966165666, 0.0087986932141379, 
    0.102502189772632, -0.418266605627436, 0.0190102707348362, 
    -0.123760132548889, 0.0904313354595698, -0.217373712024165, 
    0.102588348221313, -0.0120531243889327, -0.0103736590777774, 
    -0.0661312329113407, 0.189346973507563, 0.00347750288253751, 
    -0.0191580442379924, 0.172580026196034, -0.23526948993761, 
    0.122187225040942, 0.555118097186364, 0.156925251661589, 
    -0.286029975343791, 0.741083131271821, 0.417203506419955, 
    0.238927887985192, -0.253162655418968, 0.619943858475881, 
    0.404621440900565, 0.0045084095937368, 0.0967576002455643, 
    0.651246112982025, 0.227147287750208, 0.0383308178851967, 
    -0.00890293114430263, -0.160084119100954, 0.138665837319796, 
    0.398435325637685, 0.276209209986837, 0.111688254482802, 
    -0.0543896799345363, 0.0510817096715413, 0.00310517624276957, 
    -0.0853231838779234, -0.0913242130289105, -0.204298555100913, 
    -0.0306980127660237, -0.14390555558036, -0.14939496920839, 
    0.0253387989377527, -0.0215815733349623, 0.0362426142815837, 
    0.00274529920545887, 0.0101420034274901, 0.0122952491066202, 
    0.0102698599917869, 0.0184690053785192, 0.0216706887164098, 
    0.0692567280010649, -0.00317865887382355, 0.17201296022823, 
    0.0699547337811945, 0.133389781020785, 0.339948960613612, 
    0.210901542733908, 0.129478543730775, 0.124238860165211, 
    -0.0342400681548102, 0.632317304887633, 0.305637616978321, 
    0.0525189977882998, 0.349300837401734, 0.478107078766663, 
    0.0201125596166298, 0.757718254138114, 0.666771338243981, 
    0.051049410147094, -0.230754410213842, 1.07984365133726, 
    0.884018661510177, 0.25462114534188, 0.288921158588913, 
    0.475401283287592, -0.0165687415513817, 0.00188735956622708, 
    -0.0270505753431759, 0.564793649005505, -0.184427468084233, 
    -0.288059468842283, -0.0555081600204982, -0.194180110666906, 
    -0.136808313837618, -0.124188779168583, -0.186600589433634, 
    -0.0966899853140584, -0.187483393517334, -0.14439254192901, 
    -0.0406955072490993, -0.153140882831378, 0.0969085354205594, 
    -0.117138380616859, 0.199220739375341, 0.324042818027065, 
    0.00219348809516816, -0.0104160487294136, -0.0758686320957539, 
    0.551207713579661, 0.109638315752908, 0.163611507229199, 
    -0.284964329145879, 0.402767588541895, 0.313096974838781, 
    0.083448725257208, 0.558618679117941, 0.197528315081027, 
    -0.148530017523228, -0.212612363945549, 0.0765322829981962, 
    0.420767425681912, -0.0565952000228678, -0.0990610296619336, 
    -0.0673853228870158, -0.0756194396584538, -0.0926114393300321, 
    -0.0490848623166917, -0.0921502002460397, -0.0350587643109596, 
    -0.0822248799999509, 0.00948802183004321, -0.109873145773035, 
    0.0312885575706436, 0.0971421838776453, 0.144079724305285, 
    0.157579491444812, 0.192496995264712, 0.237219305912381, 
    0.205849503062744, 0.150946409281107, 0.174532949044563, 
    0.242986043043226, 0.237333096586348, 0.190445414398022, 
    0.166966411243812, 0.190500089693834, 0.206820321079084, 
    0.162865561811012, 0.142033645736146, 0.223398650391845, 
    0.228196983883004, 0.112853293683721, -0.00717275237423121, 
    0.286798296315054, 0.377241167546076, 0.152647732365274, 
    -0.0510162019895759, 0.479096531982843, 0.274415905737669, 
    0.011946076966342, 0.0521119320656109, 0.424919732387464, 
    0.23679210932371, 0.256194758136774, 0.897699547955678, 
    0.330149059602176, 0.127048518017143, 0.141848521669575, 
    -0.383731957526967, 0.442631222243378, 0.702564456534329, 
    0.199225405302758, -0.0771834844462621, 0.450683348608207, 
    0.338021855103928, -0.155452950220049, -0.175369383286862, 
    -0.164726005216717, 0.234553114971875, 0.23397598439993, 
    0.491327720577372, -0.00154484806340052, -0.266002263268698, 
    -0.013467390324431, -0.264183077972177, -0.0735073526119772, 
    -0.313128385833143, -0.174205913572859, -0.0910904219247267, 
    -0.209039667191108, 0.0332513014478915, -0.248332578375984, 
    -0.00211895148198653, 0.0500540139665393, 0.0528608825797704, 
    0.052509350804715, 0.0671066559746109, 0.0647250034329323, 
    0.0101171255555218, 0.0590871002771083, 0.196792453358611, 
    0.25194257949342, -0.107273876270505, 0.579948270830241, 
    0.322516707243372, 0.0586644646089351, -0.303358636776194, 
    0.0016794405186608, 0.647546591949415, 0.0915452562693729, 
    -0.123237007427928, 0.114272011585428, 0.434508249873298, 
    0.0444843414501764, 0.108095097760485, -0.165195512365503, 
    0.29287000606372, 0.180610091339668, 0.00284970681503026, 
    0.199521705813935, 0.273368461968307, -0.0307797686406858, 
    -0.115111505309651, 0.0116579366819359, -0.140324846918422, 
    -0.0170900932665072, -0.0933241390707001, -0.0237264506306201, 
    -0.153172698520816, -0.0672727590952745, 0.118641211776791, 
    -0.191497753516844, 0.180403761419221, 0.107657928426896, 
    0.0287867301464657, -0.0670986930783951, 0.321387703887337, 
    0.194839800716091, 0.060373676631513, 0.331084113391604, 
    0.123689086442744, 0.0278734337618443, -0.356252326019332, 
    0.822761497729306, 0.3016452552268, -0.0429192165360896, 
    0.229057895139357, 0.76760280231661, 0.439738050633763, 
    0.373467440687618, -0.313056613721623, 0.3933538820292, 
    0.329398934401852, -0.0242224030840506, -0.10979756050503, 
    -0.123277988960552, -0.106940587721242, -0.128730795545046, 
    -0.0965596045384109, -0.0787474939481642, -0.0488032767745635, 
    -0.126265888756486, 0.0461599600653998, 0.0301366114148926, 
    0.0767861888110235, 0.0332670141552828, 0.0614201641748181, 
    0.0368074972436015, 0.0543073701405875, 0.0270343986095879, 
    0.0720956183787288, 0.0338213450054361, 0.0815167075265391, 
    0.0655211044561699, 0.0730513349437626, 0.0766651813235086, 
    0.0806461874333227, 0.0763334883931496, 0.0851093157815573, 
    0.0907026631529107, 0.0891995616854833, -0.0446110729560783, 
    0.293092636656694, 0.213502008515842, -0.0191973536791096, 
    0.0389630634826007, 0.373078452374562, 0.263935352668683, 
    0.201674333525659, 0.304547204513837, 0.277886779511711, 
    0.102716103244023, -0.301393251509972, -0.108314414331837, 
    0.813252569813934, 0.098403583781232, 0.0117252552568915, 
    0.172791678047685, 0.0819939154067097, 0.0932890630897532, 
    0.591114859040001, 0.0980043410411711, -0.0834088989896103, 
    -0.283794046393037, 0.112524359486506, -0.0714490214978331, 
    0.119100199555245, -0.117570419324114, 0.117641471888352, 
    -0.110082437937431, 0.15282632300768, -0.24325553527075, 
    0.142430830964016, -0.0351495422204425, -0.0112996613391043, 
    0.0298453885576905, 0.0951414176982227, 0.030314978836674, 
    0.0119527241610454, 0.120126283278035, 0.101183598345893, 
    0.00641506533218861, 0.091653387054587, 0.117805929292908, 
    0.099675863455783, 0.108308317912044, 0.149406147498122, 
    0.130173336027759, 0.0893679152186488, 0.139052412521087, 
    0.174784440761738, 0.112971668458589, 0.0346995557307127, 
    -0.0363835067857657, 0.0517706056522641, 0.0388627594334987, 
    0.0551834709982814, 0.0611828214639647, -0.0199015788950385, 
    -0.00967820709265521, 0.0632085790998481, 0.148404556062155,
  -0.0826893545738525, 0.421733842165734, 0.501389526284099, 
    0.115086701863828, 0.0139255638801098, -0.214213439312611, 
    0.490704721312675, 0.386455521723013, 0.104634432214993, 
    -0.213475248493167, 0.0079139617895613, 0.423142392372185, 
    0.175862766123769, 0.0799988476586649, 0.0672866024299031, 
    0.51604975393456, 0.0478217269976368, -0.0787540187716838, 
    0.243007656617524, 0.361505352421823, -0.204299847708299, 
    -0.083188046918069, -0.0871137303548087, -0.0643981704669999, 
    -0.132250368974331, -0.164853190061646, -0.0827129677847612, 
    -0.100899231136202, -0.133056236597855, -0.156088790658126, 
    -0.000903351386874904, -0.144581942424062, 0.0255587864663958, 
    -0.0457395181672935, 0.0364538524835977, -0.189977381208422, 
    -0.00931071623702449, -0.0455635796800384, -0.000158182370982335, 
    -0.214911011899264, -0.0574843216334215, 0.0871195423337514, 
    0.041736801321986, -0.0294123839882199, 0.191727303537488, 
    0.0857496283530774, -0.0333991351158941, 0.0365230653248122, 
    -0.119485821321624, 0.345215558168135, 0.492061852289368, 
    0.00574456561731462, 0.41291143819374, 0.581866178331213, 
    0.133033705299801, -0.338273086122551, 0.296643248844806, 
    0.304990294547908, 0.301194938813685, 1.0084532506648, 0.332063899665641, 
    -0.191121025288095, -0.156669413719261, -0.395337736802585, 
    0.204037455350349, 0.51810956123755, 0.283372601979067, 
    0.105687800198735, 0.536046392655496, 0.0667605512261129, 
    -0.162886134448621, -0.120687522501753, 0.00711257501110749, 
    -0.261414149776095, 0.0363836255414657, -0.0782766670304164, 
    0.0939421317864979, -0.0440722857045231, -0.235250913569065, 
    -0.145192580385872, -0.0218974361101099, -0.115663666607449, 
    0.0211242618017913, -0.136359821327753, 0.00328792591415693, 
    -0.129257370858443, -0.00676219086332237, -0.0927330282768249, 
    0.0110266609570045, -0.103518239784508, -0.00694530932549521, 
    0.0588162133211347, 0.0733202117121725, 0.0887961305329604, 
    0.113785878270267, 0.0856784276599604, 0.0364203050506721, 
    0.088014051904078, 0.232166815528684, 0.088249924634421, 
    -0.0109197513500287, -0.247342187090211, 0.501365135050292, 
    0.514478982374901, 0.186531435313578, -0.242545826290845, 
    0.220106567352136, 0.336956681816135, 0.175294923583735, 
    0.743878742240049, 0.380778754227118, -0.025393640166482, 
    0.210260272238424, 0.640977067310513, -0.151193255926354, 
    -0.486738643605039, 0.181156994518098, 0.471849036767916, 
    -0.119738448883275, 0.0571718231052506, -0.177254406559212, 
    -0.198855199404199, 0.102705697963519, -0.169037630153519, 
    0.124293531389497, -0.160132465390347, 0.0759177640052561, 
    -0.107778780957045, 0.0864360023399583, -0.243569941339727, 
    -0.0096977076686928, 0.144896096992836, 0.224436131093636, 
    0.146495904675468, -0.00763693118681288, 0.169347507441464, 
    0.496257902306448, 0.371156378421854, 0.172571093404414, 
    0.0581927882225125, 0.0880428747410393, 0.29775241325702, 
    0.421296030305297, 0.402744302945284, 0.346220906173634, 
    0.328372012778241, 0.39624389708126, 0.363484949084054, 
    0.196038168437069, 0.183158619516271, 0.49001627412789, 
    0.349029917037121, 0.0958179713609049, 0.0673655716486618, 
    0.496009992502966, 0.212116053096067, -0.0798956092103669, 
    0.183129807627745, 0.524756720692687, 0.0437997325214218, 
    -0.190763933908629, -0.0758446587893928, 0.516422838875008, 
    0.34352179952792, 0.117820917412096, -0.212950992711458, 
    0.0374777476748879, 0.395309268795461, 0.26670117280958, 
    0.222978808173915, 0.271015277651315, 0.0972461415490286, 
    0.0124629366289023, -0.00688214959795148, -0.0406828288020178, 
    0.0950112600250177, 0.0173430278198939, 0.280321545906161, 
    0.132063099617902, -0.116767269715316, -0.200408622294717, 
    0.0847663200928585, -0.12830569310922, 0.0814400292037445, 
    -0.11427106625797, 0.0926794009344658, -0.333247530151786, 
    -0.00814156855276123, -0.178904039592708, -0.158626041702059, 
    0.0100989803834843, -0.0377806010269038, 0.166493029135006, 
    0.264855554563034, 0.0821440638916337, -0.0584289962220177, 
    -0.121623928268876, 0.25539817006668, 0.434841267002263, 
    0.230859887683325, -0.244234078230652, 0.21445588122535, 
    0.498812984335885, 0.434272600925519, 0.373526055562393, 
    -0.133451632970286, 0.707561775996937, 0.335535779267003, 
    0.0678677708808423, -0.239147974951135, -0.0431296712596075, 
    0.699948983968762, 0.221292714543441, -0.0387321529660639, 
    0.0805648539317063, -0.516014131306184, 0.262007516111913, 
    0.342149115942612, 0.415094164565018, 0.640196311324403, 
    0.159869953517116, 0.0202126203662385, 0.390828592963329, 
    0.137635087904359, -0.111929965631323, 0.250773074127838, 
    0.170780409760449, -0.0988149391799652, -0.0663144470562417, 
    0.35146080787976, 0.16417172635244, 0.0734329999067326, 
    0.0591988637722666, 0.0657406624455738, 0.0937334279960926, 
    0.0734769717239701, 0.027913115759351, 0.159226786337685, 
    0.0401974081957368, -0.0153216324163845, 0.0543218789917586, 
    -0.0694213846794471, -0.0179724744683294, 0.250869517065917, 
    0.448111680396224, 0.509292225335369, 0.265755048709699, 
    -0.0813669868803091, 0.416827664148715, 0.355979067567279, 
    -0.00881491741595457, 0.054052466751165, -0.281882480662107, 
    0.985436689486921, 0.0402859099670065, -0.093237314939141, 
    0.0483453476909183, 0.20730462214443, 0.385310585821961, 
    0.757327534333504, 0.194364773274097, -0.0623035078023332, 
    0.0308154513252809, -0.127163043745132, 0.162809500344415, 
    0.110141925216589, -0.00765858789363746, -0.0427567779635073, 
    -0.0729729917647703, 0.116646374640085, 0.0874183934668858, 
    0.0152517043932426, 0.181940553070798, 0.199005637284092, 
    0.00244233008429962, -0.119495820573088, 0.0334882432896311, 
    0.131329938467146, 0.022760275435704, 0.0569224882687532, 
    -0.158877316969709, -0.0162258979066073, -0.106853577458805, 
    -0.0949950494933932, 0.0161145685383548, -0.0923237104015912, 
    0.0514035752869406, -0.0488070289403948, 0.0781378797542133, 
    -0.0756532760207326, 0.0682268527456094, 0.0699412015186836, 
    0.0785635749272282, 0.0703185316111956, 0.0740118155105105, 
    0.0661291440419172, 0.0773311116189888, 0.0948896514357317, 
    0.0819471839323507, 0.0205561878531823, 0.074836797092137, 
    0.186358557782495, 0.137114721717537, 0.0134183558144185, 
    0.271496611025897, 0.213361593693391, 0.117827949000952, 
    0.211804220583457, -0.00491817228473768, 0.249467818049359, 
    0.524526765938586, 0.123845973294114, 0.532567576069873, 
    0.458264825509562, 0.190575794948633, 0.749410604271684, 
    0.350247605004239, -0.117186034393694, -0.0522469989247912, 
    -0.103923981646493, 0.350607563830539, 0.0238867177851596, 
    -0.07478316314728, -0.0342730144600009, -0.143429051073942, 
    0.0331911885464333, -0.175620697109702, -0.0514975306441049, 
    -0.104903266697453, 0.119113653648963, -0.0139226923588913, 
    0.127048321100515, -0.181027093969508, 0.00470065370197825, 
    -0.0392562848393223, 0.0351408281675648, -0.195470249500859, 
    -0.00728884141546649, -0.350449966851595, -0.177678129009054, 
    0.0063469424610257, 0.0366980522186725, 0.0714952663687002, 
    0.129358310337573, 0.135232793663682, 0.106941324511083, 
    0.133885323793145, 0.191246862786268, 0.144317814631502, 
    0.0871146155325033, 0.171697883709636, 0.178625289228946, 
    0.174851090545554, 0.310993522025485, 0.336201247744832, 
    0.176056500656482, 0.149858407321095, 0.473070772951069, 
    0.361265499539535, 0.11292644860686,
  0.0900303543783018, 0.126452927506083, 0.155621247457575, 
    0.174569752874733, 0.157160776100384, 0.146883716508451, 
    0.238327022998792, 0.251326935840778, 0.124404944547011, 
    -0.0426069892906822, 0.44326893267174, 0.257650575852363, 
    -0.0441102183316403, 0.0545575892123859, 0.479054924172952, 
    0.360759013624909, 0.268982466970524, 0.221044233392627, 
    -0.134400471076331, 0.518157550216516, 0.330329030381575, 
    0.0842129399321375, 0.124480058634881, -0.252989682891183, 
    0.293356173638099, 0.249731876746405, 0.469079998857782, 
    0.409556986556077, -0.196847604243775, -0.0896251323042864, 
    -0.252175117657713, -0.0186661607786065, -0.262650038093015, 
    -0.10689167390392, -0.201371613790979, -0.147517719094864, 
    -0.137193631102189, -0.155998832143941, 0.0143385793393724, 
    -0.21438209239829, 0.0938023205383838, 0.021727387136184, 
    0.0682168444315169, 0.0452977076502784, 0.0742548476173532, 
    -0.00120809321271798, 0.0594361893071566, 0.0330306563653565, 
    0.0617653447432005, -0.0389138502212855, 0.0390840506858904, 
    0.0909920730982705, 0.0834473175759376, 0.136803244683405, 
    0.157473847527775, 0.0595914386639197, 0.154063235339174, 
    0.284276402226838, 0.147751163731626, 0.168268841143988, 
    -0.258226800853225, 0.174177339579688, 0.374573029346457, 
    0.433855171117294, 0.312119368883412, -0.149951005590025, 
    0.469383566842386, 0.379402049705027, 0.107135341549915, 
    0.27200903006995, 0.384890056614018, -0.00172669555246628, 
    -0.1297861133044, -0.0714814476435039, 0.197522280675351, 
    0.435187725974679, 0.0195329534649293, -0.12229301384998, 
    0.0241050630469913, 0.27157955844371, -0.3516270408276, 
    0.271714902633409, -0.36658108346951, 0.0425732716500206, 
    -0.361302568489035, -0.118672812995349, -0.0456877902169804, 
    -0.0782113811068749, 0.300770595672214, -0.258750772270042, 
    0.0576988192448451, 0.106224514646772, 0.0604136332062021, 
    0.117723073767618, 0.166339617713258, 0.123660605394155, 
    0.111290604344102, 0.162346080608093, 0.156470080658112, 
    0.11138591827365, 0.156663477879638, 0.165235295333685, 
    0.148659292453931, 0.19651596442072, 0.269603811570762, 0.20862181062703, 
    0.109752767598345, 0.176895892243994, 0.327297294611087, 
    0.288924988761127, 0.177648476883968, -0.0753514660744899, 
    0.26739896031638, 0.340296207868795, 0.102992781735726, 
    0.395367913908384, 0.535271022862337, 0.290092027888926, 
    0.241541930439282, -0.441577109974496, 0.394381215530818, 
    0.512922216671308, 0.107509748456667, -0.0708209640866675, 
    -0.130108248117752, 0.354763728904847, 0.184521733340949, 
    0.656330733778452, 0.891907755622228, 0.0608217687610491, 
    -0.124815092156487, -0.06639028915676, -0.0193644404330411, 
    0.035739782359042, -0.0273574331342213, -0.0683562320504845, 
    -0.0565507743438315, 0.139368094447219, -0.112513354189653, 
    -0.0490947651646294, -0.0455536964675697, 0.055107365616801, 
    -0.130313399268886, -0.00436617601182086, -0.0653888569950606, 
    -0.0796220054634078, 0.0223878348188319, -0.019820179068969, 
    0.0934617374934806, -0.104179350108571, 0.157380028300609, 
    0.169253738892956, -0.0459083403745065, 0.354455479135931, 
    0.210074825553245, 0.0241012351942552, -0.0416776142417847, 
    0.0825223645086918, 0.600522939007185, 0.0203728604261325, 
    -0.178350127663025, -0.0215308643187675, 0.305463053374154, 
    0.0464762343802514, 1.32171422216653, 0.612055814481901, 
    0.0439916205456595, -0.323246340746537, 0.509214786413433, 
    0.431310328493916, -0.447153180490154, -0.185495334540334, 
    -0.0115363474920815, 0.118220188121401, 0.0380647513734106, 
    -0.00335651537284434, -0.000706804038724834, 0.00405074638715701, 
    0.16989547713372, -0.119956136362539, -0.084455427165124, 
    -0.0176343396692728, -0.0510736030998926, 0.0329034777457715, 
    -0.0982145533165469, -0.0642033024377166, -0.0181896860026245, 
    -0.0574635529441523, 0.0294324303094955, -0.0758192488131322, 
    -0.0303215806401736, 0.119671339133573, 0.138861840660447, 
    0.106541553598471, 0.116647363084107, 0.124231134182602, 
    0.0998461835333296, 0.108811593038442, 0.109925200917211, 
    0.0974926371122218, 0.17523979085576, 0.189154875733083, 
    0.167918786423071, 0.190426126082433, 0.203376776932763, 
    0.168078939332737, 0.236133094083971, 0.286728459510045, 
    0.135821600621331, 0.0585501742311307, 0.560601319306477, 
    0.127253347904296, -0.151284648499089, -0.173074647918279, 
    0.534312981401637, 0.44823695309016, 0.280342503016437, 
    0.462331939572489, 0.499015772169915, 0.25337212851084, 
    0.131691913927629, 0.70325052747447, -0.0669998751733632, 
    -0.232269766081415, 0.327174160062905, -0.0621607560262733, 
    0.629940352260467, 0.0143635397711305, -0.0439473217034914, 
    0.338750926513898, 0.148548629383243, 0.145624191070432, 
    -0.0438897571143702, 0.211338725065886, -0.0403282142437888, 
    0.17792245692934, -0.376860127335213, 0.0309782420046337, 
    -0.341566380683843, -0.240415829220118, 0.0115997371712734, 
    0.0889298323222394, 0.146679152738865, 0.188752486945477, 
    0.267796725255439, 0.334230795000745, 0.263974446962879, 
    0.175194680214479, 0.259947960280323, 0.36728936932629, 
    0.281451071332392, 0.202542742371438, 0.172525129784135, 
    0.172548134571262, 0.129113404648142, 0.109995999690684, 
    0.108781834714248, 0.171286678103891, 0.186175703351075, 
    0.127831962638218, 0.13269077863649, 0.129408808614183, 
    0.123564341365402, 0.258236169022912, 0.221450731826859, 
    0.038679785391279, 0.341690557649739, 0.358710422974337, 
    -0.141193471157387, 0.0194441979479872, -0.125861302094337, 
    -0.264372422651492, 0.630847103052112, 0.347114464121481, 
    -0.133485575806108, 0.131225703116012, 0.81842051396438, 
    0.367764304891443, 0.0542672004124883, 0.462676659633913, 
    0.486548970240078, 0.174473474505453, -0.0118859703717384, 
    -0.0311333523711576, -0.176781723210283, 0.0902306917565108, 
    -0.0375200690958185, -0.193517082847151, -0.0465965500741584, 
    -0.0901205440830442, 0.0777171239939886, -0.141008883398807, 
    0.130169968574774, -0.0464701721629221, 0.115902255736061, 
    -0.175578065390677, 0.036723572457058, -0.0771452633227877, 
    0.0258439388055647, -0.228091921026848, -0.037912731197379, 
    0.0596900932778597, 0.116482337435306, 0.140418291033125, 
    0.147143855973324, 0.150853369435349, 0.170233436735836, 
    0.16906012387913, 0.129395752540541, 0.114909013399917, 
    0.203577850903365, 0.217332097496671, 0.190911772395066, 
    0.213592074099958, 0.25382010150984, 0.232472691529903, 0.21726871462452, 
    0.209359314154027, 0.14002771412403, 0.211169477253165, 
    0.415657664232046, 0.228498979374026, 0.0200448283870743, 
    0.445463657141724, 0.333887657628595, 0.0510183873492663, 
    -0.0964581690954845, 0.580725793049096, 0.327956262195326, 
    -0.00904574787758071, -0.0644281932353938, 0.0811104233112336, 
    -0.312750745106566, 0.390352516966264, 0.504911944347675, 
    0.250876719622809, -0.354921744702566, 0.414500575742562, 
    0.298841532549711, -0.036067053356097, -0.212528942399549, 
    0.115924191674322, -0.343135558978758, -0.0201829148102107, 
    -0.272509748809094, -0.161277964970213, -0.130297389598416, 
    -0.19828964007001, -0.0354727304241079, -0.191535776726516, 
    -0.00875201386997321, 0.0880232129543, 0.109375614952995, 
    0.129519902639472, 0.147632300529602, 0.121935919531341, 
    0.0804081697223122, 0.114927671190871, 0.0999041515351799, 
    0.0582865244186555,
  -0.0189362911035373, 0.131382788303818, 0.16014157658536, 
    0.113268686330399, 0.0649875659300965, 0.0687893238956772, 
    0.151201845033746, 0.150580114322927, 0.109081730928139, 
    0.0725532340870558, 0.0883136755520633, 0.138580897740247, 
    0.151674851901538, 0.114898576328522, 0.0952197390647497, 
    0.146402827893078, 0.151385899069383, 0.13333912092355, 
    0.148964666595769, 0.132535954107575, 0.0442210595429982, 
    0.0221841699571459, 0.0664012443447476, 0.0201958918108759, 
    0.041647367547913, 0.017246484732268, 0.050458026515107, 
    0.0254847185665085, 0.0729646454315308, -0.0207367162185933, 
    0.0493307238141454, 0.137771768130358, 0.169326128783237, 
    0.10068790728826, -0.000976084820820677, 0.249542711193461, 
    0.197101712121999, 0.0312225946528738, 0.199151445738254, 
    0.514527513501525, 0.314229769097744, -0.11158663886627, 
    -0.303874068534832, 0.727607543145972, 0.574151335810369, 
    0.102528380978304, 0.118097093749112, -0.0931490953891538, 
    0.787048936977843, -0.0483369152560231, -0.127349837830102, 
    -0.320819554622226, 0.0240866032370385, -0.0687485632949945, 
    -0.0261880825503623, 0.0560186790663751, -0.139012187511843, 
    -0.0923861629278514, -0.128061375488219, -0.0419420446374538, 
    -0.156208201163698, -0.160279240086773, -0.0227644736461275, 
    -0.080526950216549, -0.300452839496656, -0.062241258555794, 
    0.00753160800275843, -0.196997072205696, 0.411804752387269, 
    -0.297207225487571, -0.00258404182165024, -0.0672061271931837, 
    -0.064987908788406, -0.0194979384063702, -0.0387072184611498, 
    -0.0374602110209545, -0.133085877352126, 0.0913430552915372, 
    0.226908947193482, -0.318498663076646, 0.257572105090579, 
    0.686792637863001, 0.129401231852072, -0.195720567424859, 
    -0.00425475381931241, 0.575947017597071, 0.274460162737853, 
    0.17253775793663, -0.25635074040539, 0.28263198160816, 0.36614273165794, 
    0.185320691282246, 0.109346250639983, 0.184146826542406, 
    0.254891221924671, 0.171228901535339, 0.0902725888898036, 
    0.114801530635294, 0.207376667610945, 0.144626370942196, 
    0.0354152365530815, 0.0261156570215388, 0.0390155841864083, 
    0.0337117182569376, 0.0385999846170068, 0.0323628764322524, 
    0.0393558274600688, 0.0362687696276703, 0.0415670352919632, 
    0.00850570934050627, 0.0852758372599471, 0.0655084703990676, 
    0.169900216772336, 0.264882940062916, 0.169602040941036, 
    0.0802470396454943, 0.307169657899868, 0.292621193381251, 
    -0.0111891520657286, 0.408241362612604, 0.719142375001406, 
    -0.252107130748934, 0.383476757340994, 1.03812961250681, 
    0.012120438068021, -0.532659583501301, 0.269218547269117, 
    0.522763217026619, 0.406728667240467, 0.932332021254555, 
    0.493247476202492, 0.024526166749033, -0.00820664597030178, 
    0.169155943439766, -0.281401148431394, 0.611562651634825, 
    0.178156716999904, -0.207331923698602, 0.239657738993818, 
    0.45501389147958, -0.0484740459863869, -0.0301137411520879, 
    0.0240377346440926, -0.0653958588377747, 0.0424598847657289, 
    0.00245893179616943, -0.0174293675240881, 0.0593160116625346, 
    0.0132296181975534, -0.185410931252695, -0.0887877946866366, 
    0.47345636784679, 0.211791762121687, -0.188015303145994, 
    0.198237896099455, 0.318339991412564, 0.124879553348339, 
    0.544271183805956, 0.334374068043689, -0.00509824243469836, 
    -0.137403400931673, 0.0312695613688258, -0.239764735818336, 
    -0.117370796749016, 0.0332548754028143, -0.123646682775845, 
    0.0852149575622225, -0.0956197315936204, 0.0657506723864821, 
    -0.0729798265931679, 0.0988948835700818, 0.00406387855765536, 
    0.0330578920520683, 0.0436713919119328, 0.0520869203260534, 
    -0.01077239464538, 0.0326572147284549, 0.0398966049246282, 
    0.0333095115069069, -0.0567378188587057, 0.019111249209145, 
    0.0669716663648542, 0.0541778272488123, 0.0547917416922505, 
    0.0887937029832478, 0.0846265307907336, 0.0979010350237496, 
    0.0954417565905948, 0.034768964714989, -0.0947291735339088, 
    0.390508861396528, 0.320948280431846, 0.189711390903085, 
    -0.165757556540623, 0.224530007371163, 0.351103102162145, 
    0.228728592544223, 0.463030713287814, 0.306771443669394, 
    -0.220695737850431, -0.0114719720077722, 0.581662341817806, 
    0.298055615836843, 0.0921986124125594, 0.27242132328553, 
    0.501216067222704, -0.174335769146335, 0.33997115499206, 
    1.03525140248192, 0.05812933653496, -0.128672566756079, 
    -0.0582470770946085, -0.0190109582666155, -0.0912173673056902, 
    -0.121533728642401, -0.16059167108681, -0.154516653244332, 
    0.0274065002662775, -0.0673196085125673, -0.0236005266778991, 
    -0.139715934990815, 0.0207364970202294, -0.1903350856888, 
    -0.126552262225048, 0.0685947724875581, -0.1028756083216, 
    0.0811206703442238, -0.0519215149665995, 0.0654930701296247, 
    -0.145770085900891, -0.0124211364788573, 0.0498779557579751, 
    0.086173828280643, 0.0404012234652573, 0.0294567942868855, 
    0.213522753055587, 0.0788757479445011, 0.153465239385415, 
    0.323973014015722, -0.0782831427572626, 0.74202820044957, 
    0.482154550311737, 0.177391120752148, 0.100613039650419, 
    0.259910071938488, -0.249397075616678, 1.03396355275259, 
    0.351583295267824, -0.32354276219213, -0.283530023415927, 
    -0.525909721276318, 0.53303067196569, 0.34686794932229, 0.12314500683455, 
    0.047039993667235, -0.0697314321079208, 0.248392048094879, 
    0.954054825704475, 0.11615186285885, -0.10839357317659, 
    -0.155407268763761, -0.155011220663022, -0.11118304769684, 
    -0.129025340615352, -0.134655748553168, -0.115592587522155, 
    -0.115643553389052, -0.0580752947954454, -0.0657350377574082, 
    0.0583364218916118, -0.301642290796378, 0.366086695400842, 
    0.231897066466604, 0.0594797854975612, 0.0396159122592603, 
    -0.223835869743566, 0.189252134313119, 0.497341614452768, 
    0.317656257113962, 0.0954090043487755, 0.0241122131773501, 
    -0.356103255567649, 0.726644574752301, 0.391703854250611, 
    -0.157085735515814, 0.831548474047339, 0.302418572855328, 
    -0.127683153138093, -0.0759416530219301, 0.281940141740059, 
    -0.271184306932347, 0.116791721222438, -0.304980379372151, 
    0.105213713812186, -0.312445055602205, 0.0285659687217898, 
    -0.383446693011985, -0.155143545772504, -0.112529050325724, 
    -0.259201598086876, -0.0344124524113777, 0.106073426756972, 
    0.198064046134339, 0.209866770216216, 0.216457586758431, 
    0.21279125413944, 0.177714583785951, 0.169823063784116, 
    0.269519344224374, 0.291259832663536, 0.174003950551904, 
    0.13095628145421, 0.10946402430951, 0.111641576734281, 0.110068185793277, 
    0.11415021691487, 0.10684440434249, 0.108261336032113, 
    0.0770234270230838, 0.0733773150739768, 0.0845343989258928, 
    0.0958372279112481, 0.0980604176074529, 0.10628014683902, 
    0.120012645451353, 0.0934377754916309, 0.0887091713938502, 
    0.17075850610577, 0.0875040300530894, 0.00282116313877483, 
    -0.0207707554344101, 0.000477116139319014, 0.626969571262445, 
    -0.0130550380047106, -0.250124892242976, 0.171838892762062, 
    0.412592875835163, 0.0746327967454521, 0.241874563371666, 
    -0.2390927578906, 0.360072760586334, 0.48210293282493, 0.262360641081679, 
    0.0107819212074907, 0.337915578149587, 0.671949608781015, 
    -0.132745327191173, 0.706375734705305, 1.14103605016871, 
    -0.0215358052862375, -0.144046275521718, -0.114302768951341, 
    0.0519642566504372, -0.122302631253602, -0.0962755755169903, 
    -0.0745447219378058, -0.0237281885317635, -0.158226414496534, 
    -0.0343364909354194, -0.155010038547517,
  -0.208219384033128, 0.105416448612095, 0.67387824258865, 
    -0.024721191842311, -0.215052945303511, -0.0711857715176822, 
    0.62455433928111, 0.200309734826059, 0.114814370230665, 
    -0.133018348401842, 0.292750814593579, 0.335053772860792, 
    0.290730108206447, 0.124814788464006, -0.0914813251338261, 
    -0.140555942419473, 0.510193380318276, 0.161304626852016, 
    0.0466066759826195, 0.216345515323266, 0.0984629665303879, 
    -0.149904156616183, -0.0499957803458533, -0.109249324360664, 
    0.0671710658901778, -0.0185396224356494, -0.144891851961302, 
    -0.178088358897358, -0.00436162504523038, -0.110158431059221, 
    0.079599458991288, -0.105878107333115, 0.111571626548709, 
    -0.0906220608814638, 0.0672008989465424, -0.12168655821444, 
    0.0153170579346279, -0.0668307021059889, 0.0287082438956488, 
    -0.199199594910654, -0.0168289055443878, 0.057724534918119, 
    0.0827936230997415, 0.0773066975949858, 0.0826634960654018, 
    0.0555132435074963, 0.0320148247362748, 0.0936236045137311, 
    0.0907145000778927, 0.0109209374177204, 0.0731254287149402, 
    0.136646329347085, 0.215483482094783, 0.314455547511336, 
    0.198339178562725, -0.00245396661651034, 0.390335346307113, 
    0.272907795458852, -0.0838216466952199, 0.0911352312371601, 
    0.604828966091759, 0.208876566794942, 0.171906964654973, 
    -0.253833368967009, 0.833572201426274, 0.590605746056989, 
    -0.253143455310734, 0.722519308770027, 0.649894882069711, 
    -0.112135792675265, -0.16666304488106, 0.0852514756075135, 
    -0.104558412458232, 0.0933340000865549, 0.0380277300840062, 
    -0.118152310532963, 0.141746961825996, -0.016361219550404, 
    -0.123052478708134, 0.145614070763276, -0.0291257890436934, 
    0.161142913546816, -0.116690236494689, 0.10241352571832, 
    -0.369034643427283, -0.0689661286806006, -0.114633906849219, 
    -0.213520997891774, 0.0463879688427079, -0.201551090993744, 
    -0.0327764961365231, 0.0456497400635675, 0.0158077809390479, 
    0.0166885637516345, 0.05598928677855, 0.0296985188018121, 
    0.0420576698303569, 0.0503613613701887, 0.0447470168054868, 
    -0.0121060345564676, 0.228941926698609, 0.156604796376041, 
    -0.020694178302535, 0.296831735307667, 0.247080805750321, 
    0.233994158361667, 0.457646999876753, 0.165344834558273, 
    0.00736475488873939, -0.142545641005549, 0.313365118240781, 
    0.499357866150759, -0.315362189909212, 0.0836400672569918, 
    0.793878174724815, 0.45177420440344, 0.0508429656535069, 
    0.711916358633618, 0.851359239084416, -0.0146907621633943, 
    -0.170670085107823, -0.0909245525825753, -0.122853130988758, 
    0.0264017074208304, 0.0746642347108342, -0.00767562188510337, 
    -0.187900759334653, -0.309865185748825, 0.0387873565670039, 
    -0.168743278288867, 0.0631259734626762, -0.143104266919294, 
    0.129592294918688, -0.103630781412158, 0.13284161646475, 
    -0.114240273556708, 0.11607576018342, -0.0991825163019988, 
    0.101517813858498, -0.21357057084436, -0.00097394350585546, 
    0.0547040061511476, -0.00727037184731419, 0.0477022891438715, 
    0.127376572973188, 0.119129190784319, 0.122782835892789, 
    0.112066221758855, -0.14831386654174, 0.322912774508337, 
    0.462280995971426, 0.191667855244866, -0.428374234343077, 
    0.128730293184052, 0.519795886339633, -0.00323204259014005, 
    0.240731368289339, 0.898197154336072, 0.389765325195408, 
    0.224907865439492, -0.0685251984626017, 0.407649598307237, 
    0.270831502031946, 0.227759282893866, 0.194811773870257, 
    0.0652997390675171, 0.344329894559479, 0.214474084093153, 
    0.124358952661847, 0.41981018437818, 0.204623276394566, 
    0.0615540859777657, 0.0320539889593933, 0.0287376697069534, 
    0.0280753146431996, 0.0484278021559496, 0.0620657071570133, 
    -0.100607235258463, 0.103893368254679, 0.158298537234963, 
    0.139805670307654, -0.126881051639704, 0.117392933367313, 
    0.471855536092085, 0.385672697432387, 0.18220527958981, 
    0.0440119459748778, 0.344151553625589, -0.175749202576929, 
    0.360354356629735, 0.734771753504242, 0.102923139447986, 
    0.0274116015551924, -0.0916694095581351, 0.391094233245217, 
    0.225319360987612, 0.278701038374797, 0.696099360151473, 
    -0.0268065759053435, -0.0579276467763234, -0.225842296701439, 
    -0.100147904016545, 0.00455141443719644, -0.139004751686757, 
    0.0903312631870642, -0.144269350363583, 0.003470121456394, 
    -0.101086857111583, 0.0205062765626358, -0.187085022086865, 
    0.118771462241501, -0.0426162732437838, 0.419285822976098, 
    0.294584118412076, 0.116298341461809, -0.265898782174389, 
    0.227631151601219, 0.445203759411675, 0.212163747050343, 
    0.0903963911231449, 0.0206445869301548, -0.0215733475104389, 
    0.276248106339872, 0.361153923515127, 0.189076826207756, 
    0.367343352097049, 0.752943127727179, 0.4761298588379, 0.145793673636924, 
    0.0751903816811175, 0.594095323749985, 0.491071154760641, 
    0.145534537287693, -0.0654473015452758, 0.239483759250834, 
    0.44209296405723, 0.271673057265826, 0.0971013177925826, 
    -0.230808020139991, 0.0550838820386466, 0.589587844341557, 
    0.051492025506882, -0.214819856597237, 0.111222824560443, 
    0.428427051769265, 0.073430128737679, -0.323158457520392, 
    0.291142794608978, 0.625389114517136, 0.140555221761752, 
    -0.113316984268189, 0.146908747769749, 0.11606865256397, 
    0.0340342102118842, 0.141638547232031, 0.0625087708959722, 
    0.126127816416892, 0.179166539712224, -0.0315232686984012, 
    -0.0164519250309943, 0.0751060247424045, -0.133199813355219, 
    0.241500382943551, -0.246463851596077, 0.141959793341131, 
    -0.381524966997766, 0.0428181163155326, -0.23731684372927, 
    0.0737642998052055, -0.405183647310212, -0.00305059813154125, 
    0.0196564528975678, 0.0366258179755917, 0.227161891974626, 
    0.252461502362357, 0.126382106666816, 0.0423154233259861, 
    0.135547714895585, 0.233334236768937, 0.225506486650974, 0.2908638404366, 
    0.298480297444853, 0.271536897672139, 0.280502657705054, 
    0.322326041443588, 0.291373583248222, 0.231870809884634, 
    0.260203792081203, 0.349098761109091, 0.321539817430148, 
    0.162610710356726, 0.135690381845614, 0.679169936778985, 
    0.329499439541867, -0.035020212788226, 0.355652924675576, 
    0.472949869905047, 0.0669705793617427, -0.0136825309198333, 
    -0.148916439484378, 0.464422777215519, 0.815450458331258, 
    0.269601367478561, -0.00226992366596029, 0.382384028336639, 
    0.314186981884292, -0.0235032521514831, 0.169957964307165, 
    0.44189727032912, 0.0189442685455378, -0.0393876670614721, 
    -0.0155815953072663, -0.0159031199884053, -0.019653584908808, 
    -0.0172924355418581, -0.00274394222253285, -0.0285940851428673, 
    0.00702617310312514, -0.0129736245430926, 0.0591162784014436, 
    0.195865749004151, -0.0738494337776283, 0.0363200769876127, 
    0.444083739299808, 0.207741373499648, 0.0374242852220777, 
    -0.0742393489049066, -0.0856433364484179, 0.330697911163092, 
    0.328956110618471, 0.412317508253099, 0.247575961497204, 
    -0.076507610663151, -0.119693424786897, 0.328760061483663, 
    0.414141844525669, 0.209917941540752, 0.246598231826712, 
    0.557402735897557, 0.108584990634512, -0.0685961685010617, 
    0.0188729062336875, -0.169157944302488, -0.0133935279861987, 
    -0.0812865949299272, -0.00639572269061592, -0.224523569109872, 
    -0.0828715615373246, -0.088161409407735, -0.295007667533369, 
    0.0810787018058854, 0.147775527392554, -0.0280450651527135, 
    0.101588290681529, 0.410753984201348, 0.156299538888526, 
    -0.0628928888601813, 0.0806047944928779, 0.495372493790281, 
    0.0909586273059637,
  0.00120425158679131, 0.0663990176757441, 0.0617035538632768, 
    0.0792112935238045, 0.114097608037812, 0.0951052612134455, 
    0.0889740574894752, 0.124931069729992, 0.100392282840272, 
    0.0848742036139405, 0.169090418962513, 0.0344405167977394, 
    0.107118106031139, 0.465617084522931, 0.23701959915599, 
    0.0393840059531911, 0.0569332548959451, 0.580995962931753, 
    0.00886394661220297, -0.0947818360924873, -0.0526682127000338, 
    0.439432512163984, 0.176832659982288, 0.121280752062767, 
    0.646709133488385, 0.353917723829815, 0.193198373331372, 
    -0.0708651911758882, 0.600813785984661, 0.187103445213876, 
    -0.0425471849589887, -0.0427771875794587, 0.0676201865162389, 
    0.0733145632013167, 0.0223729169309361, -0.0823627098214635, 
    0.287715766552824, 0.134913115772858, 0.000885816589422772, 
    -0.00831984411323668, -0.068252689901882, -0.118230516440469, 
    0.066028227946961, -0.22642035405596, 0.0312054441842073, 
    -0.240161581399044, -0.0792490384500961, -0.0628532338059396, 
    0.0737688397732158, -0.267144395557378, 0.0630637784989783, 
    0.0651912592939263, 0.0537246945455405, 0.0945698298544617, 
    0.125029491733207, 0.0892466997962728, 0.040796024637425, 
    0.0684445369618385, 0.102122048498898, 0.0462783331243595, 
    0.0955364389568701, 0.110658812651481, 0.122984208013694, 
    0.161118880974224, 0.192411497491721, 0.159754151287387, 
    0.107899167209196, 0.143180313742486, 0.226746245367833, 
    0.239749620884998, 0.175539950516307, -0.13015471138723, 
    0.16324072183518, 0.46058044604216, 0.241293015123848, 0.069542352030257, 
    -0.0400732299615172, -0.138698024197695, 0.566411650616575, 
    0.165861961821805, -0.0343063916995205, -0.170142172051647, 
    0.274108257242371, 0.382065562802142, 0.602758687405939, 
    0.462691673201957, 0.00286021650032453, 0.211090106789272, 
    0.876733644527054, -0.0385113715602426, -0.146236472088322, 
    -0.0440761098322548, -0.14043653527733, -0.0443180642200383, 
    -0.135585543800408, -0.111829156467877, -0.0984934748313331, 
    -0.0701263839107086, -0.181392270637742, -0.052756761091352, 
    -0.0656124867469937, -0.0117301538872622, 0.0378781797897367, 
    -0.0113485650390025, 0.0825133643689333, -0.00187054790862484, 
    0.0487770961831619, -0.0375946936239945, 0.029791261541043, 
    -0.0285023957537384, 0.0601272173814013, 0.0189403782131685, 
    0.0797590752765377, 0.206654376504251, 0.122085540976497, 
    0.0590715381598903, 0.272096166192029, 0.225412757760064, 
    0.132492883937209, -0.429207690694559, -0.0480175844469508, 
    0.631608004194841, 0.349635230392538, -0.128265052020237, 
    0.0499003328812941, 1.18500293447938, 0.385008367139631, 
    0.516290697456745, 0.357500477340092, -0.441659630963565, 
    -0.392237180612375, 0.0213620404026822, -0.148146179954918, 
    -0.122385122736584, -0.0888913515655758, -0.178164689056516, 
    -0.128101302943622, -0.0472116545369808, -0.237066804826636, 
    -0.0986457654369532, -0.0950516908174809, -0.063843033893181, 
    0.133724815111945, -0.130588196217251, 0.108655123034746, 
    0.00503369516277428, 0.0567284137384147, -0.0320222416836116, 
    0.0220820621632954, -0.161533046504704, -0.0556569497312985, 
    0.0553794290827904, -0.00344093116270573, 0.021576311245643, 
    0.0386915594095533, 0.115288918648955, 0.0353863181502338, 
    0.195144939240913, 0.271197315370389, -0.177155670796797, 
    0.2343349310402, 0.406100770075149, 0.54832713904817, 0.563958593938567, 
    0.246155767372544, 0.5533209291472, 0.730880751050414, 
    -0.224841320368847, 0.781143029785904, 0.873173975186961, 
    -0.254153510354152, -0.112046088982087, -0.1150253369008, 
    -0.108102978737282, -0.140182859685944, -0.0813291423857686, 
    -0.0873497930234041, -0.0556018238402484, -0.0494234736162499, 
    -0.0315033244305369, -0.0233417420289624, 0.0797037523616111, 
    -0.115580467249559, 0.0567590877182649, -0.0943247339117616, 
    0.0329437064475851, -0.260070220009553, -0.0672680036328884, 
    -0.010023857543237, -0.198502003200769, -0.0167488544572002, 
    0.0359868406386617, 0.0680525320891437, 0.0617985684321569, 
    0.0551844897529496, 0.0558834857280765, 0.068317749384689, 
    0.0830922900036088, 0.0631143732476125, 0.0406901307266217, 
    0.155624055751209, 0.111730957487382, 0.185960815953092, 
    0.175323236356801, 0.187944191729233, 0.469195246792887, 
    0.28478815941724, 0.010146922380806, 0.356884480747518, 
    0.317473845438254, 0.184687035970915, 0.816802705419816, 
    0.354703697052237, 0.193648442925592, 0.528450832462443, 
    -0.0316290438775079, 0.612095803415145, 0.558729919856857, 
    0.230172079895769, -0.0866770671322563, -0.34784391255033, 
    -0.198129236049198, -0.0478138957195074, -0.241062792332901, 
    0.0426662231806283, -0.216077591460522, 0.0533994356948028, 
    -0.0970497171481498, 0.113613940987321, -0.226517384172352, 
    -0.0289973536277717, 0.154884545874428, 0.202978132290106, 
    0.14198196098566, 0.153000945556534, 0.160655886576875, 
    0.110012647661429, 0.0883314071557218, 0.206710591563217, 
    0.221140711629977, 0.18558615874743, 0.171553475290543, 
    0.163083865564858, 0.15450575363451, 0.145589397542403, 
    0.144935564526905, 0.166058945911602, 0.1941741094679, 0.172411883036757, 
    0.14172987774881, 0.176850794748196, 0.166465062386009, 
    0.118893231375789, 0.219685304552919, 0.291186133009115, 
    0.154225765003286, 0.087131226967106, 0.326347148603791, 
    0.362224437832463, 0.216469840959355, -0.127682860269129, 
    0.547127869230384, 0.275591251540087, 0.00728964903202868, 
    -0.128406331575614, 0.438280258095674, 0.43866520614386, 
    0.421644647688331, 0.200849401074118, -0.277202447575132, 
    -0.106761360904601, 0.524194212978721, 0.456399838685508, 
    0.231785544148257, 0.0976117060311276, -0.00080772940144494, 
    0.674993469796383, 0.110487346835004, 0.112061741423386, 
    0.312757147335976, -0.0151452584585079, 0.148951968422637, 
    -0.241311206084914, 0.049407739140993, -0.394353253801066, 
    -0.15366683204375, -0.0536009684455631, -0.206680425835656, 
    0.101306227562455, -0.297256800348931, -0.0323142653487255, 
    0.0917998765610098, 0.117484619650716, 0.139783777513232, 
    0.262366953980742, 0.257407890371533, 0.136061624866352, 
    0.0570667936730657, 0.199690441254928, 0.416814018869264, 
    0.2424731033976, -0.0509501384954926, 0.0144904882725751, 
    0.523435771699055, 0.357392032971602, 0.119182049426846, 
    -0.130214106779918, 0.0471310414247758, 0.51160454767965, 
    0.287100730234975, 0.149929540625048, 0.531664405200837, 
    0.281532842293969, -0.00205426752029247, -0.0671588921951282, 
    0.614464755085586, 0.296734966391531, 0.117040158228876, 
    -0.233629581406536, 0.241703101128975, 0.487471813221159, 
    0.116351920884379, -0.116383899024382, -0.0212461264306102, 
    0.372960307366287, 0.325006982184737, 0.252167958762393, 
    0.180873930057036, -0.205643094531038, 0.267108624068579, 
    0.384490458953549, 0.180603376402511, 0.0654260466669551, 
    -0.032501344123046, -0.22583740907642, 0.276746898802775, 
    0.531775959557831, -0.221877902042386, -0.227741760034545, 
    -0.0561585778646585, -0.0990231323121871, -0.189959762519529, 
    0.00178493479272544, -0.221490202621762, -0.0235210673117033, 
    -0.169448096412159, -0.00480967636582633, -0.191060950559944, 
    0.0280313459138752, -0.0971384577256202, 0.0832222414501334, 
    -0.0725193691517375, 0.0180293986407258, -0.060995553703714, 
    -0.0234936987577925, -0.00298988515443144, 0.0280671638845126, 
    0.00912891207529486, 0.040017309368784, -0.120315608841992,
  -0.458589359205646, 0.108758273365038, -0.287891679006723, 
    -0.0378538855385942, -0.33977740666163, -0.129090007572045, 
    -0.233277906786188, -0.245799445531332, -0.0283133778440013, 
    -0.243130988362472, 0.00381600967137894, 0.0750816953144428, 
    0.0617978633455919, 0.0831614908242187, 0.0672435268925879, 
    0.09150421224534, 0.0758004809000111, 0.112690293217795, 
    0.0838935967840745, -0.0435499707245633, 0.25557988126164, 
    0.0104726546489044, 0.52536835309875, 0.546487343820759, 
    0.0550371690762524, -0.250403336071708, 0.0656440897132582, 
    0.656467814092069, 0.278753289366279, 0.0871027237376098, 
    0.278647650006736, 0.224068346280926, -0.289324252406741, 
    0.247414510673604, 0.701385008564341, 0.193619082652582, 
    0.013563857124298, 0.320273298773981, 0.177233576325339, 
    -0.141778211187664, -0.242754387958674, -0.109639879268893, 
    -0.189621353162405, -0.166996536777186, -0.0363803542641765, 
    -0.1865065718893, 0.0456678090456722, -0.101220976985702, 
    0.110195871990593, -0.184797064601684, 0.0955002968934996, 
    0.0871004403759664, 0.0402559590497677, 0.161759806036378, 
    0.201821892835902, -0.0414132000248884, 0.310235337328603, 
    0.427575247955649, 0.173570314024473, -0.0228004891677275, 
    0.324182193298355, 0.901428040683442, 0.199153116808668, 
    0.0728697671229583, 0.0882506082365135, 0.131231695239665, 
    -0.246233326357814, -0.0409382476369645, 0.213804345011126, 
    1.04624955299737, 0.918201982680484, 0.283499020454765, 
    0.0606063757721797, 0.0582499421444495, -0.206514950957847, 
    -0.0036574324673195, 0.157274816010361, 0.233830095345503, 
    0.519504608098085, 0.0331630198849484, -0.228821796613724, 
    -0.0890503921505768, -0.0875333409760411, -0.107249824154182, 
    -0.0879114371317868, -0.0263366467300733, -0.12618407609725, 
    -0.00348133294618883, -0.0970374874925194, 0.0238819845626269, 
    -0.0737925652502464, 0.467485651436942, 0.226705828458164, 
    0.240753500215457, -0.294387954002945, 0.487362181423954, 
    0.347377807611628, 0.0321274431634112, 0.0756169876294367, 
    0.502255479292279, 0.297572085329119, 0.138702542559006, 
    0.0840708308799164, -0.0574719838280124, 0.414047520434067, 
    0.0746142017415273, -0.0998040349502532, 0.137050873352106, 
    0.277763583375783, -0.0399922147011622, -0.0732360441133876, 
    -0.226876858181171, 0.102636564304352, -0.166102459595431, 
    0.0360679106791883, -0.230595534834843, -0.00459287733089757, 
    -0.108246356285059, 0.0604754154844308, -0.320878993825929, 
    0.0273392705268435, -0.0724698973240032, -0.034230896251914, 
    -0.045790195930113, -0.0424674857193559, -0.0846034577527316, 
    -0.0394470874229904, -0.021251414246124, -0.120923793835367, 
    -0.224839061523908, -0.167614220062955, 0.950728737825035, 
    0.0456807693343104, -0.195688084243709, -0.41899310139857, 
    -0.0911079204758004, 0.696250805595846, 0.531295575942213, 
    0.579140391028759, 0.679534977932898, 0.00339782712485046, 
    -0.061814984704547, -0.0939920988377925, -0.0152447274105445, 
    -0.0692174921279467, 0.0129565609430209, -0.108402591081255, 
    -0.00505070565832265, -0.0681506118736218, -0.10944177980952, 
    0.0949925321108193, 0.00447820881782088, 0.0964943045290322, 
    0.00211460895331968, 0.0326153902114044, 0.0182599899925516, 
    0.0171859993484247, 0.0868831375302197, 0.0409278745151544, 
    -0.00406261963664389, -0.159345261664407, 0.046610936593272, 
    0.334011276606042, 0.17965224167696, 0.072189587117578, 
    0.374707489073488, 0.257458486608875, 0.0224493638447101, 
    0.368385787625065, 0.306954396966581, -0.0941660547737716, 
    0.555897000981462, 0.505300930999499, 0.0879127072908985, 
    0.515098053135996, 0.608065567773913, 0.107774300578306, 
    0.0839530802641588, 0.780908077320033, 0.161537773877528, 
    -0.0285302989434605, -0.00236818383189227, 0.00413239593326387, 
    -0.00669958084525606, 0.0028276015079514, -0.00272156310128878, 
    0.00136680092589517, 0.0109745349273502, 0.0441390543836905, 
    -0.0137723220222007, 0.145454420905658, 0.021573839611585, 
    0.26731764126102, 0.26931430748542, 0.0628534074567794, 
    -0.0197548888825596, 0.421781655340832, 0.267379639495367, 
    -0.0647586663993437, -0.146551768279422, -0.0791104797655795, 
    0.658745977609118, -0.0235905483475618, -0.0821821257775312, 
    0.196420725447586, 0.377643477292222, 0.0100807784542588, 
    0.931568123613121, 0.525495612877074, 0.0379779476333208, 
    -0.139531669514786, 0.0617557262557696, -0.0838180795931503, 
    0.0156567330715559, -0.0817202210676277, 0.0135134582938338, 
    -0.182055807759031, -0.0579159741298247, -0.0207209039926458, 
    -0.217767027967798, 0.0417282617778433, 0.206553415879579, 
    0.13983519367089, 0.00972533953442284, 0.104011826834808, 
    0.325566986801006, 0.353761458535697, 0.345265987225594, 
    0.291441128575273, 0.158702492929197, 0.0689733939348394, 
    0.108915560645875, 0.558561439930387, 0.635693946143502, 
    0.324689055864627, 0.131591661045054, -0.276274740492363, 
    0.618840112923437, 0.56690882513704, 0.0141825638593156, 
    -0.134703756183573, 0.0216444918171586, 0.690283313668201, 
    -0.0812732006005935, 0.0203287465676808, -0.186550248344596, 
    0.147813919401921, 0.500018930394974, 0.266479979102654, 
    0.0944195371624921, -0.191977476701894, 0.38440169162352, 
    0.243123907136042, 0.218887645715595, 0.246581955242496, 
    -0.220238781420411, 0.293971818183548, 0.37948683994206, 
    0.0858430843983722, -0.122381399108497, 0.311964144740958, 
    0.422484342502276, 0.0242825916870722, -0.0521136314204598, 
    -0.115104847920259, 0.18854287212583, 0.271538532133351, 
    0.0976415578394226, -0.0407777829588778, 0.140671061120785, 
    0.072236514149553, -0.0801595971083336, -0.0719374022971138, 
    -0.0408159808027151, 0.030119439010643, 0.0612575796997372, 
    -0.171514036468373, -0.079412346821118, -0.0743361801106547, 
    -0.096106080099819, -0.0519252155989669, -0.210449775006292, 
    0.00460769953408877, -0.168942918124523, -0.0122717819560574, 
    -0.2497291237528, 0.00785617235931194, -0.122845585241805, 
    0.0106516124525768, -0.245976296763847, -0.0274880600067377, 
    0.0639459616058301, 0.0632416235473841, 0.110708690966351, 
    0.157384185013936, 0.127629912481242, 0.126664344383665, 
    0.190122403569411, 0.167845844515131, 0.115955274876179, 
    0.169592679646308, 0.18008402248577, 0.254902836127771, 
    0.302396130543658, 0.206195049519569, 0.193335919034156, 
    0.377359987503012, 0.244489843076188, 0.0257581418732976, 
    0.279881482781596, 0.454068201492244, 0.322239816597562, 
    0.428915304385415, 0.373652903602653, -0.0505050945956205, 
    0.636510134419258, 0.467354356108664, 0.141433729668091, 
    -0.0979925108203095, 0.382679486401355, 0.298767635508528, 
    0.247086281404709, 0.248263779583104, 0.0381668330321619, 
    -0.110185085859768, -0.0859416634776018, 0.305715173704778, 
    0.108554831565975, -0.053065673301472, 0.160241401039316, 
    0.258082361052033, 0.136367411533098, 0.0726887695789796, 
    0.0563735074949442, 0.0531745032296904, 0.0547838986946611, 
    0.076176810535886, 0.0664911708889961, 0.0494395799512643, 
    -0.128733852330198, 0.35374146298734, 0.217056109922456, 
    0.00649841426797718, 0.234473224799805, 0.214694636115277, 
    0.148368764818751, 0.574203709159327, 0.425862047797737, 
    0.0458839540065844, -0.370551028705567, -0.0137056588060286, 
    0.584696766086978, 0.257390702237315, 0.118943589469489, 
    0.952845485957157, 0.282348212354678, -0.139029986131098, 
    -0.481673117723121, 0.264875476208909, 0.563906395452041,
  0.113746994426998, 0.229411971771142, 0.141673427478994, 
    0.0647208530803271, 0.0283358739275607, -0.0495799991225684, 
    0.30843880108239, 0.444909008404374, 0.0335914796709518, 
    -0.123282884020163, -0.145802567617622, 0.363971257005486, 
    0.37283833664058, 0.343114029781118, 0.182183257623714, 
    -0.18948558209856, -0.133412893586969, 0.639127705777785, 
    0.408101848066412, 0.106597137462244, -0.272858919685624, 
    0.0134788182858554, 0.509133184609595, 0.0912550907165126, 
    -0.00587264652072937, -0.0404708731638629, 0.51902922283522, 
    0.14096957092472, 0.0961761532541668, -0.165636079654262, 
    0.0902599725946931, 0.44095571011916, 0.0669253096555388, 
    -0.0781333780366785, -0.136719059958196, 0.420528992366933, 
    0.125429310042396, -0.0607824127985015, 0.0595176381197739, 
    0.275880057694668, 0.160076901535392, 0.219496926969477, 
    0.13811493679028, 0.0237192757077803, 0.113503081988472, 
    -0.0242214898526085, -0.0889138749782012, -0.122118283080052, 
    0.00798856824427086, 0.0983251021938003, -0.0428642294438944, 
    0.0198769440826475, -0.0281612961991819, 0.0373539549048665, 
    -0.109497824995019, -0.00297082243498784, -0.0527845480507613, 
    -0.0355433822600113, 0.0935204930194232, -0.0951554054974704, 
    -0.143735441355294, 0.247022643411418, 0.193020076568036, 
    -0.0194819650588371, 0.0347570516991214, 0.369201208444583, 
    0.310336851749759, 0.13263012519621, 0.126152485172113, 
    -0.0951041851832517, 0.821134196396956, 0.130190123297097, 
    -0.521607669207131, 0.209974970376482, 0.683185125487931, 
    0.800617360801635, 0.517954004655531, 0.00797341207033142, 
    -0.404388375639887, -0.119089643216224, 0.56550533219516, 
    0.762821495292805, 0.352620925190098, 0.0470362546798568, 
    0.0396548382391027, 0.24579468138658, 0.371723974138153, 
    0.25074151227208, 0.120585168603092, 0.0991437648318556, 
    0.219080673306912, 0.229088876177067, -0.0654553613480345, 
    0.00336635678526535, -0.152919384518254, 0.184911030401898, 
    -0.0522810570528628, 0.0504597795163826, 0.0173502720331852, 
    -0.0240238690336202, 0.0326264735598226, 0.0230242524204575, 
    0.0809456033191572, 0.137397817262827, 0.126449781008403, 
    0.0727516957639951, 0.0799605342850131, 0.212451398053336, 
    0.0797370168519827, -0.00763448546165128, 0.17127105956674, 
    -0.164938060418972, 0.27636672124784, 0.507942136620502, 
    0.0412611753798088, 0.0205764489361094, -0.102975065642207, 
    0.576273759544084, 0.123482193540341, 0.0819194081931772, 
    -0.231304775429381, 0.162044880552689, 0.448699866357765, 
    0.0322813270227045, -0.0547022087695203, -0.113081398449649, 
    -0.182043332911672, 0.352052639686727, 0.39691593562774, 
    0.190391954359117, 0.110819021391708, 0.294794186698466, 
    -0.0525193823611853, 0.204098739632224, -0.166138341414953, 
    0.136920927936305, -0.146406500161155, 0.094400596125488, 
    -0.273603937921851, -0.0672049313168866, 0.00168771418701257, 
    0.102509561373927, 0.047312838668884, 0.040824683375468, 
    0.107203435704971, 0.0761279065252051, 0.101070469349573, 
    0.0785284095555231, 0.0749434767563382, 0.00104171113392042, 
    0.0365506374208219, 0.0993310588826419, 0.0737146136538051, 
    0.091161717043235, 0.189953103899624, 0.11630168550452, 
    0.0204848821177454, 0.272991920860182, 0.249697643729062, 
    -0.234811356200277, 0.0381153724450475, 0.44957889424838, 
    0.584625887971472, 0.303775949231654, -0.247498513514329, 
    0.4142844427415, 0.373701950059109, 0.202299656638629, 0.622135509434788, 
    0.136846683229287, -0.227201960554897, -0.159059280519552, 
    -0.0159255975294701, 0.0709593610921657, -0.0161099869466104, 
    -0.00681495682568525, 0.158746924314243, -0.00402616689836592, 
    -0.0921475931997536, -0.121920550055268, -0.363194596859746, 
    -0.129068284398579, 0.109864508029962, -0.289626762976407, 
    0.189049729841681, -0.116883703306786, 0.0169986398653595, 
    -0.0122950292264104, 0.085997625414587, -0.0951549793652516, 
    0.132844890253645, -0.234292011593785, -0.00761373176278245, 
    -0.126111889923204, -0.0426651072237844, -0.0828751376277586, 
    0.015861337483262, 0.00347086460659242, 0.0934344750440354, 
    -0.0818713218464844, 0.0798097423631956, 0.0637977945823462, 
    0.183586479435086, 0.10667433760188, 0.0317722333136226, 
    -0.038507416184544, 0.161179992418364, 0.111722128998742, 
    0.0407942473090506, 0.0158430342475923, 0.0663140117665073, 
    0.177842538943397, 0.355965520186376, 0.00538005874402774, 
    0.133275143941542, 0.873580139180862, -0.00248816926420206, 
    -0.135575842275472, -0.108036790887119, 0.675699790889437, 
    0.195222094719328, 0.0125178571673943, -0.228068942169976, 
    0.0663908502765502, 0.657735231662721, 0.671537912688394, 
    0.24426976401833, -0.344362565570666, 0.342602647084124, 
    0.43631536654532, 0.0202607961646904, -0.0346143907970366, 
    0.32151969270902, -0.219815966846408, 0.0115041585847645, 
    0.499576445693668, 0.274915197734554, 0.113946647755553, 
    -0.119484888613432, 0.127143774642193, 0.218076605408312, 
    0.131359278920107, 0.0888354018312415, 0.0785915917934457, 
    0.0785696234956702, 0.0796466425234232, 0.0860895533515501, 
    0.0822673699610072, 0.0469532774832974, -0.00672146636963075, 
    0.26470656531074, 0.167930807584766, 0.0604106356544693, 
    0.111883994875437, 0.535368856828045, 0.56321871013713, 0.08821629974563, 
    -0.168698548894692, 0.113879493370686, -0.184401717744336, 
    0.68655996022821, 0.540491017193242, -0.0527183300319314, 
    -0.0804378498366137, -0.0655361516813264, 0.712277458607752, 
    0.122291866044865, 0.194755110855371, -0.122847534609069, 
    0.348179432901904, 0.276314752454482, 0.136047423903186, 
    0.0785940881275737, 0.0712113598538889, 0.106176951747238, 
    0.0965036711474776, 0.0539376828672791, 0.152411293761398, 
    0.0856313734118024, 0.0273646844461819, 0.0690536315224249, 
    -0.0471402235826701, -0.0320051698143399, 0.513830851382051, 
    0.313308797660639, 0.0583716751463654, 0.10650651384682, 
    0.648373005528351, 0.104530594886197, 0.00440051794247429, 
    -0.0137744563936829, 0.365043351180012, 0.500687510171153, 
    -0.000523397996585587, -0.181508588747112, 0.456047821474852, 
    -0.409425597475419, 0.827774180412498, 0.363924471958475, 
    -0.0878781149302877, -0.262154796513404, 0.156773759508634, 
    -0.217766828262392, 0.0708188255351129, -0.409875047289428, 
    -0.0174274014429707, -0.358307300155967, -0.139191322700468, 
    -0.209206237471722, -0.11674462423131, -0.0404934982101023, 
    0.166465344163484, 0.0134066480419166, 0.0316427332879092, 
    0.0790235521094374, 0.121769925194811, 0.10272189963777, 
    0.0919928514494233, -0.0527666885125616, 0.0360210404892787, 
    0.0241431936781035, 0.0428229848714499, 0.0537713300495549, 
    0.0563875299903266, 0.0512982376704004, 0.0601663829962782, 
    0.0382213762573505, 0.0818022551098971, 0.0529863339305165, 
    -0.00417976084442175, 0.252387303356439, 0.148340046035837, 
    -0.0604611859109975, 0.493318678647928, 0.304480452214289, 
    0.0760136586236957, -0.0282661682859965, -0.267343600526975, 
    0.157147694561723, 0.71960264850885, 0.205842803101664, 0.45014710264886, 
    -0.615937260846371, 0.725146201469196, 0.336632120521984, 
    0.109303944850418, 0.185950654844107, 0.0126706695368473, 
    -0.156400390160826, 0.999046114892786, 0.456676247940103, 
    0.0625995444135912, -0.00913863401546658, -0.0181069233250503, 
    -0.0193016513680985, -0.0270779914699355, -0.0309735694158771, 
    0.0406424041063835, 0.0217472710347474, -0.10854895928974,
  -0.00586945690815198, -0.123141809486036, 0.0520407302685404, 
    -0.0563705647719284, 0.155723190922213, -0.259097835848081, 
    0.0872135913254636, -0.153722370448932, 0.0428036953721858, 
    -0.314650729494754, -0.0581987230527196, 0.0052524849955753, 
    0.0630478334627037, 0.072744000737057, 0.0578538292981971, 
    0.0367162140264134, 0.0527849502985413, 0.120100532744284, 
    0.0847783727678045, 0.022810144205758, 0.132324640896626, 
    0.139568113055143, 0.168573362365989, 0.278818209816354, 
    0.255755675966846, 0.181563798731645, 0.377353831868659, 
    0.425876137446757, 0.149838273855612, -0.195742435027873, 
    0.282225140724282, 0.45761675853023, 0.449477546773962, 
    0.467953234553902, 0.0971893249160473, -0.150902990732868, 
    -0.287790796472112, 0.533157620050479, 0.411322193144894, 
    0.183502006130528, 0.115300714742741, 0.220946086852265, 
    0.11365502419618, 0.0497722068893871, 0.035268759666865, 
    0.0322036581097902, 0.0306783849247029, 0.0283000215408192, 
    0.0193809703830905, 0.00375837344068185, 0.0763333079652968, 
    0.0966420016742602, 0.106107675443178, 0.115021723185696, 
    0.119841104179572, 0.108211485806496, 0.112694778302812, 
    0.141525870162147, 0.116197105367087, 0.0759897705823645, 
    0.181600276476993, 0.175735010419225, 0.0828371245274143, 
    0.203459738765584, 0.324589949456676, 0.202700718266502, 
    0.310355714349074, 0.325881124655576, -0.0797789602203925, 
    0.23880902266502, 0.669742175504122, 0.0698583360751976, 
    -0.173960680644462, 0.350806550077963, 0.271597568862542, 
    -0.106581204494198, -0.279108530358895, 0.132134268326168, 
    0.357536801343841, -0.0650399988973584, -0.101816918318402, 
    -0.146712018036007, -0.0185197858355682, -0.162333793329303, 
    0.0103593941888449, -0.15053019988519, 0.0266524440851751, 
    -0.133857177632035, 0.0521562169931346, -0.139288347578485, 
    0.0717618161337307, 0.0643970000504993, 0.076775873877788, 
    0.106045541272405, 0.11203792883273, 0.0728764510570698, 
    0.0917380096554514, 0.106774990539299, 0.102104676847414, 
    0.048005750824997, 0.0781110179122006, 0.0962979132263647, 
    0.106209082298777, 0.140315602646893, 0.160114541171622, 
    0.108578482551251, 0.0488624545570889, 0.144176265753208, 
    0.273850137850147, 0.219835716112084, 0.00348070782666496, 
    0.509420140823895, 0.269701743151601, 0.066380867316139, 
    -0.152252181343597, -0.00738072864704344, 0.594018574953629, 
    0.2807010175687, -0.0202977610003708, 0.266344486187027, 
    0.292042621177564, 0.156031133632013, 0.129387790016203, 
    0.262024093142238, 0.491172203678188, 0.255330702029775, 
    0.024025412330997, 0.211607169201304, 0.278061019088322, 
    -0.0318678245835942, -0.0265192424411277, -0.248989918781683, 
    0.0850884224490643, -0.0959994284621486, 0.0593103084510264, 
    -0.160047563553947, 0.0980722471980495, -0.213791802130142, 
    0.078901360049777, -0.227911371659716, 0.110560198041081, 
    -0.0628740958825711, 0.146597060034698, 0.321502463764658, 
    0.149993859597816, 0.0173543787760687, 0.0724003265779387, 
    0.311888921243043, 0.0129113397777304, 0.141370047227609, 
    0.84273431820899, 0.195666233825175, -0.1001090968043, 0.232871217776954, 
    0.900881610516939, -0.0136689577290901, 0.206873020837677, 
    -0.221266440024969, 0.701868463489695, 0.335178857578981, 
    0.259856479715048, 0.210538220298959, -0.386817515550399, 
    0.022344631348758, 0.691680771023795, 0.173173176057632, 
    0.0632027932064362, 0.11115415736944, 0.320354442532865, 
    0.804690763663034, -0.371898569763189, -0.291530297030958, 
    -0.18399518429887, 0.51625605010999, 0.264156101157038, 
    0.102974907040636, -0.2237224986747, -0.146245245681865, 
    0.412161439584836, 0.267362391584076, 0.123236101465116, 
    0.195928046921919, 0.0415878339828811, 0.196005964972726, 
    0.361842571752431, 0.0258298230068445, -0.0511418889337972, 
    -0.00846630633826033, 0.216864074197132, 0.155769662949502, 
    0.148512952383405, -0.0988935861824364, 0.0475970168299493, 
    0.304080168785147, 0.152007002739748, -0.000190534475945275, 
    0.138263610341946, 0.223789468127857, 0.237324723506736, 
    0.164540203130863, 0.142126472904438, 0.521564430990997, 
    0.0734220693578717, -0.0114903226271338, -0.106513392520508, 
    0.33666245545927, 0.264732622029177, 0.373065331030025, 
    0.160773196956796, -0.158720535436023, -0.186249259720076, 
    -0.0420055555025303, -0.153289242376911, -0.140971480292301, 
    -0.0694712492433592, -0.159737280840122, -0.0655666005697562, 
    -0.0990682020105752, 0.0180417956342107, -0.128857213056588, 
    0.0704333000908816, 0.0271094997670238, 0.0667517844025931, 
    0.0101758879054627, 0.0605525827233707, -0.00531620619082046, 
    0.0530545487101073, 0.0209341753850849, 0.0612739216038347, 
    -0.0561630372906208, 0.0415112906574676, 0.0743698473924297, 
    0.0675098597190508, 0.118333405474121, 0.161896891972532, 
    0.124196755564216, 0.109416331728229, 0.11056672943642, 
    -0.0183685507538144, 0.229374380788717, 0.398590408318374, 
    0.130724354322305, 0.0901159248717545, -0.31888641029971, 
    0.125860597531625, 0.666846568178001, 0.175791275117217, 
    -0.257170197388316, 0.185370683160453, 0.479701541416669, 
    0.132806261900522, 0.0365068785692995, 0.104511595519107, 
    -0.144832288309581, 0.81693946909219, 0.529457608697224, 
    0.152587892057147, -0.132251837167133, 0.849145547703782, 
    0.170380620376265, -0.0229766415473941, 0.035704308264801, 
    -0.184926710395535, -0.0282907350821872, -0.0274289486253102, 
    -0.0853653409305378, -0.134229667672661, -0.0541491734277934, 
    -0.0770116990148458, -0.179114353771764, 0.0325157905345923, 
    -0.0878942518928774, 0.00283212230394959, -0.0706348471289216, 
    0.0200952364747802, -0.0662079765543652, 0.0199363774858465, 
    -0.0570343234694556, -0.0105937497049401, 0.0225845616087518, 
    -0.0469674547576335, 0.0117866890030237, 0.165318763102831, 
    0.317565578465622, 0.181934796337462, -0.117331806885737, 
    0.131264663676289, 0.439236544546175, 0.0471272543979457, 
    -0.0529401549445059, 0.208766223202024, 0.269795698355447, 
    -0.105548763509355, 0.671174164339507, 0.748067599829059, 
    0.248809335664794, -0.25388884353902, 0.289905852806109, 
    0.512652400523818, 0.359426337423878, 0.204587596525138, 
    0.0610661530142303, -0.0783732403616775, -0.0670984084888622, 
    -0.0434661807570139, -0.0690791932014436, 0.0213326850362723, 
    0.0117378259789665, -0.0967524064819198, 0.0802222096291315, 
    -0.066111534518146, 0.0421707881899805, -0.225637708502613, 
    -0.0865356450907517, 0.033494453343423, -0.125175034359537, 
    0.0626701407885335, -0.000925371579956716, 0.0933559272987618, 
    -0.0874894681322139, 0.0660108148001776, 0.0465275104291258, 
    0.0523256479809858, 0.0587384244576276, 0.0646241597585561, 
    0.0505851653208589, 0.0597132300337307, 0.0611783133070023, 
    0.0595249160077896, 0.0171288934567467, 0.0214630278554587, 
    0.162448738667051, 0.24594190149283, 0.119196559728329, 
    0.0489886897808042, 0.444641611136361, 0.135357382762535, 
    -0.124808392091642, 0.161427674753853, 0.37134737783668, 
    -0.0496652562666628, 0.403825797243263, 0.624022068393821, 
    0.293693710101363, 0.206258842305125, 0.0574351821853917, 
    -0.111846292119497, 0.419866944476373, 1.11742541611721, 
    -0.0457422893431444, -0.292991017103349, -0.00790502993874302, 
    -0.216349967385362, -0.0341630563933541, -0.222819697917041, 
    -0.107480671087298, -0.0479116474271806, -0.208160360490384, 
    -0.0375487927160102, -0.253522986837237,
  -0.414159534492074, 0.0799123425331782, -0.121365539395056, 
    0.00369815459608674, -0.299908623387808, 0.00243183173279551, 
    -0.266462003172628, -0.0168319373016162, -0.0112487418152208, 
    -0.0879097515309197, 0.0282125454815081, -0.00896777744371667, 
    -0.0142233704468124, 0.111169167469626, 0.0821335205420196, 
    0.0418973747067301, 0.0485010963067116, 0.114404627455316, 
    -0.0444786317429711, -0.100743304508064, 0.0340252320154736, 
    0.287231036264954, -0.0554438229917676, 0.548448617516714, 
    0.422283310728592, 0.0180290190010213, 0.328912077203504, 
    0.580195480723012, 0.166033831791725, -0.103089013966458, 
    0.224055668063164, 0.820054375431481, -0.0241511107178435, 
    -0.124357954446772, 0.0757934395193129, 0.700698215773216, 
    0.0265473875473891, 0.523924867797359, 0.775810371130195, 
    -0.106684540754925, -0.122288862445426, -0.135763368739792, 
    0.0236834638488764, -0.233521279848833, -0.0657840290533567, 
    -0.129603798319699, -0.110410116150381, -0.206968171848259, 
    -0.0697811627152185, -0.221708074605048, 0.105220996075039, 
    -0.0406241037584705, 0.0515119076311942, -0.0319229526556778, 
    0.0330015932165058, -0.0299789521031671, 0.0132723901788445, 
    -0.0373593334603218, -0.0329402158814374, 0.0120020117818266, 
    -0.0737565212442461, -0.0558766380204321, 0.00302506204592524, 
    0.00477519570952735, 0.0332615267742626, -0.0707302865647265, 
    0.00503801194731955, -0.0181590008068466, 0.0294272349323488, 
    -0.0808462228782944, 0.0233887295842459, 0.0623158437663229, 
    0.0738600037230224, 0.0800858791956691, 0.0824243673703151, 
    0.0678471756756717, 0.0725144698497806, 0.0926200025461939, 
    0.0795250115136313, 0.0385527074952791, 0.0929831874788369, 
    0.132766468819085, 0.13899708920786, 0.133217023287345, 
    0.133465860874139, 0.131996750345594, 0.200648917605474, 
    0.167278601008344, -0.0257920022164334, 0.124486574415215, 
    0.450388342043051, 0.154184197620072, 0.181573288681611, 
    0.765834146045913, 0.224246475648889, 0.15981801990843, 
    -0.0632816756040856, 0.636322197245969, 0.181283270093549, 
    -0.071996760881841, -0.0398382733312024, 0.541751738030613, 
    0.259592171173051, 0.035222446097885, 0.196441855798809, 
    0.44180941849329, 0.157343640109605, -0.112904196761144, 
    0.122532365083221, 0.508874655732951, 0.240992440483788, 
    0.139321803714006, 0.282635066947856, 0.303253200497575, 
    0.154664851889028, 0.0562582535596659, 0.0641811756277805, 
    0.148822899181677, 0.0573959297899082, 0.0795861104975836, 
    -0.143379271984002, 0.004996714799798, 0.276827994350822, 
    0.481753682655436, 0.262293709629631, -0.247954773238936, 
    0.302568511018148, 0.434454627758877, 0.082220910563299, 
    0.0275611349592869, -0.148008017766935, 0.381526752316156, 
    0.210688876228753, 0.0581175516146979, 0.114831334212771, 
    0.257369135368024, -0.0344946212954099, 0.352079746605143, 
    0.412654770491201, -0.0449342791386553, -0.123098476499641, 
    -0.00604100272577618, -0.0776455501662678, 0.0688101200921198, 
    -0.180009455254941, 0.0627814999566969, -0.214410395210181, 
    -0.0411030975905616, -0.125809129447111, -0.0334931092898564, 
    0.00120334576641164, -0.0304139304815933, 0.176963155308552, 
    0.232132399596502, 0.140662923952193, -0.155061202152232, 
    0.215974598519839, 0.362801374574588, -0.172147373801274, 
    -0.209349071673039, -0.123934272826686, 0.494359090872961, 
    0.410047389779102, 0.136569198260117, 0.0368802502875341, 
    -0.679963683082584, 0.249377848869905, 1.006927397807, 
    -0.692675384747744, -0.247960304241055, 0.164707773342667, 
    -0.183163455950097, 0.24336981732112, -0.0545470313116723, 
    0.124154720352857, -0.00671310483883845, 0.0108324226733621, 
    0.0519130714184731, -0.0801133983150349, 0.06328151675504, 
    -0.089195154427327, 0.159718732672267, -0.0901182608577604, 
    0.111320502138458, -0.339456151085333, -8.49564752511828e-05, 
    -0.20911686883404, -0.181215158093313, 0.0114879538464869, 
    -0.211659916169202, 0.0402699593103981, -0.00291326350394193, 
    0.0216870201270539, 0.000616446949477628, 0.0385513265269922, 
    -0.00114466633222769, 0.0383775141062922, 0.0266912697899875, 
    0.0529436306719917, -0.0161918765118046, 0.0689568094972528, 
    0.0974818589600545, 0.10159468731604, 0.178790379797632, 
    0.17471435036098, 0.0588375264360334, 0.148999067841921, 
    0.345958397654927, 0.0930781144179798, -0.045993177962126, 
    0.289227099506673, 0.196982130411046, -0.368804280286998, 
    0.456217443204266, 0.718637874086392, 0.257817941659723, 
    -0.167263906813536, 0.508126457230992, 0.372709478491691, 
    0.1339945911597, 0.345103609973371, 0.295677396581722, 
    -0.0215397595836884, -0.0570387836635565, 0.0507606933905772, 
    0.465728801479425, 0.44515779337537, -0.0184680422197699, 
    -0.165386455829171, -0.0733203852498793, -0.0820612604436192, 
    -0.280029553677843, 0.250983653744931, -0.184993323804738, 
    0.198108637418168, -0.202520492297405, 0.129597368676505, 
    -0.132624412738286, 0.122938616567702, -0.312401819785153, 
    0.00708358747636519, 0.0287276704547315, 0.039819294697387, 
    0.208807864812729, 0.142392021403361, -0.0133862348098631, 
    0.0969062043817049, 0.303342609918742, 0.0951231169995867, 
    -0.0818857915843888, 0.593489303287232, 0.171632521404024, 
    -0.419763836018006, 0.0869272090377563, 0.647573106875581, 
    0.219251943331371, 0.174892322191922, -0.35977797143695, 
    0.410943362945103, 0.431298293445354, -0.00500615062524634, 
    -0.175599208431501, 0.171839132233166, 0.285234625161733, 
    -0.00867655483956006, -0.0334844107828988, 0.00214212867559221, 
    0.28138819304843, -0.0554581293772116, -0.0553274620981279, 
    -0.186524966548524, -0.15955651650181, -0.00828919836559502, 
    -0.164185941848968, 0.00743275574692864, -0.187378515436564, 
    -0.0407583826773278, -0.103983435440483, -0.054958583904228, 
    -0.167934675670217, -0.0613002729673293, -0.0351132642859346, 
    0.274606434316021, 0.209939846397045, 0.0283723508495711, 
    -0.115416092141907, 0.456571139677485, 0.199791690407956, 
    -0.0363256249629085, 0.0655403731825253, 0.557762905796642, 
    0.293944237426993, 0.234165664399537, 0.399513362247942, 
    -0.0632231846853667, 0.9813497355893, 0.296140077703764, 
    -0.206760733779495, 0.687406526068669, 0.274057146576698, 
    -0.428493065656121, -0.151780925843612, 0.0169104024661444, 
    -0.0953325092433303, 0.0211589426106035, -0.155371461291657, 
    -0.116471737998099, -0.117090286392601, -0.0963477876753408, 
    -0.221244390291993, 0.0862995069139121, -0.105623592118848, 
    0.0379262567901458, -0.0719708104650044, 0.0592865216499598, 
    -0.0197690823469614, 0.0970438027790814, -0.109463028375261, 
    0.0304907338657989, -0.0382589547193786, -0.00344256798874407, 
    -0.147113168457028, -0.0181998352205649, -0.0627031147237958, 
    0.00332041287444548, -0.12839348133168, 0.0162552387180313, 
    -0.136227382222364, -0.026580622164776, -0.149907015519084, 
    -0.0627704694709208, 0.027991900198192, 0.0428367314514286, 
    0.0146577450143816, 0.000337228241434034, 0.144072012777552, 
    0.121480310551693, -0.109177100012895, 0.121549249978542, 
    0.171893171406725, 0.187356079902828, 0.133171012557025, 
    -0.311527717885008, 0.607120736532352, 0.451592158129051, 
    0.204384452057505, -0.112308094058811, 0.601883161749081, 
    0.368840731154322, 0.296593239106136, 0.237695482028077, 
    -0.471363774434604, 0.0802228699097263, 0.65971558982355, 
    0.185488981058998, -0.558405147909018, 0.3265267151997, 
    0.988983595898261, 0.0242774558559295, 0.00591090072252931,
  -0.0980868211272306, -0.195981015910136, -0.0477388302571613, 
    -0.230685838394262, -0.0538301061516331, -0.187027936019677, 
    -0.0318919630543932, -0.181038136321871, 0.045224800590714, 
    -0.179826479848735, 0.0781016835356591, 0.02210980482279, 
    0.0561486323091301, 0.0265320861648405, 0.0521365698625356, 
    0.0136370871525774, 0.0373949232377766, 0.0543718992367731, 
    0.0691561009114705, 0.0224365797312852, 0.166151287004194, 
    0.0354352493761281, 0.216570358957284, 0.240223231381326, 
    0.0652851671007633, 0.103717293614247, 0.348708904750497, 
    0.170622379089715, -0.0765875232682572, 0.318700784044257, 
    0.360374437220426, 0.159202887308202, 0.389146414878954, 
    -0.406809275357371, 0.244931816293717, 0.360675647019105, 
    0.36428382914899, 0.564145026471492, 0.277561170452838, 
    0.0642560554108056, -0.165834817182716, 0.0973975359699712, 
    -0.2110910689308, 0.0884124008726335, -0.24476645843526, 
    0.00560240923681113, -0.259091195309891, -0.111284754772511, 
    -0.0751298226096018, -0.197988868477513, 0.0609209020146364, 
    0.043105566925184, 0.0731282428131461, 0.132663653242112, 
    0.18341178509695, 0.0847280997982871, 0.0710119962942418, 
    0.125954231137755, 0.121400585860977, 0.0593760343001695, 
    0.0801414863144503, 0.107374726618182, 0.122667469858308, 
    0.145828282804536, 0.148637269510769, 0.115583236069232, 
    0.123855650391436, 0.199451093687331, 0.157117616804764, 
    0.0727546221410413, 0.065300460429116, 0.0699600313120516, 
    0.291979126940396, 0.399297730058968, 0.186607151466765, 
    -0.0960093428457479, 0.30629659521848, 0.493467227605073, 
    0.245587753244361, 0.0398182144776219, -0.0571809411237533, 
    -0.370462404584082, 0.374338688005998, 0.44851109012548, 
    0.218123537879111, 0.169998945754445, -0.230052314003146, 
    0.673831997779089, 0.336060120534365, 0.0366394198799297, 
    -0.273761106862291, 0.0766069737780911, -0.315119193275756, 
    -0.0350808474118758, -0.326359707969373, -0.185740170566488, 
    -0.0320339661761815, -0.248852225167512, 0.0487936274699292, 
    -0.111642360878502, 0.181696811828687, -0.0248465948033545, 
    0.0346080868607343, 0.0548917811188453, 0.101704860769553, 
    0.0300563641574407, 0.0914996419356118, 0.0434809252395101, 
    0.0463879365393915, -0.109603651886489, -0.00453422232067734, 
    -0.00477009815872063, 0.00338955966362314, 0.00545474294544236, 
    0.00598133699553949, 0.00337791939436231, -0.00233974388085503, 
    0.0290003496297812, 0.01764000068549, -0.113414543921135, 
    -0.0549921164393904, 0.434989522082873, 0.285425075455415, 
    -0.104460721651502, 0.332148742849686, 0.39941241862974, 
    -0.00896682439547999, -0.217492432546256, -0.0939134237210459, 
    0.938630547179534, 0.0959720576416224, -0.417204191305557, 
    0.261716465885435, 0.492031698895489, -0.0471834695862718, 
    -0.237605097854462, 0.0938607818237421, 0.704776086122463, 
    -0.108834569820465, -0.00216635574902388, -0.0662436828778887, 
    -0.236944939082271, 0.339949018876942, -0.439900442939403, 
    0.108555846212592, -0.262996402978529, 0.0462429774358028, 
    -0.127219186781234, 0.149596862122239, -0.36598241997427, 
    0.00469551448414696, 0.0589455770824202, 0.0925289232809301, 
    0.223599945234541, 0.275300909896829, 0.211813723264156, 
    0.253570125346905, 0.318269531384612, 0.190728093316998, 
    0.247671719617772, 0.528897138616305, 0.254569122170215, 
    -0.0227099394335321, 0.794450355912292, 0.515647393319523, 
    0.0426793913792688, -0.306890898655956, 0.039138304888981, 
    0.789373981597618, 0.126932878201546, -0.0473762670098541, 
    -0.175602289132347, 0.376103081838485, 0.250042383741734, 
    0.17784606933031, 0.565212375506681, 0.339093797645326, 0.15163599006837, 
    -0.12477618996813, 0.403245080293127, 0.190793640586006, 
    -0.0162993371921751, -0.0656228597526281, -0.0767219777487579, 
    -0.015610806572464, 0.249517145653522, 0.102837645002381, 
    0.0565555317977964, 0.117364131610934, -0.174052628558486, 
    -0.260023741238566, -0.0946114858953725, -0.0835772490422659, 
    -0.179977192225053, -0.0436812518108741, -0.165126940923888, 
    -0.0403297573921967, -0.137159339700524, 0.0382152267943005, 
    -0.137875327042918, 0.0874536837103041, -0.0105659059831832, 
    0.0333843733116727, 0.0120216275455122, 0.0387397251719593, 
    0.0276641072309929, 0.0545978363598442, 0.00643472722231675, 
    0.0359501757854384, -0.0181220218913856, -0.00614844688572705, 
    0.123035326094077, 0.143170877305969, -0.00527044618495222, 
    0.168641579986312, 0.241178592251791, 0.158807849190487, 
    0.454744446000638, -0.0167166024738422, -0.208237833044877, 
    0.0209594624333217, 0.591255172106741, -0.0118634700178491, 
    0.205493008619527, -0.338355633434297, 0.56721577529797, 
    0.423986430414174, 0.213524284007873, 0.0223887936845099, 
    0.568340637658509, 0.122252287791572, 0.00742820096139155, 
    0.0863155392272056, 0.118099131189245, 0.00485941681912339, 
    -0.0222853971324903, -0.00418230572201317, -0.0738251724575041, 
    -0.0501661605049191, 0.216551696030679, -0.0839529463704423, 
    0.164011669536788, -0.237529694503319, 0.0172606183206357, 
    -0.0936011332658546, 0.00673022816709287, -0.327675515350747, 
    -0.0603683246450024, -0.272560695393789, -0.267689438461976, 
    0.00873606226010107, 0.0461716682021981, 0.0661132340760437, 
    0.0712304664509952, 0.119337091524151, 0.0959029090854727, 
    0.0852751166255999, 0.0900234670274609, 0.0901727737105123, 
    0.080222073883613, 0.110834474692047, 0.0967063160764313, 
    0.0943439620824514, 0.0922973035204339, 0.113271240826077, 
    0.0968293490365726, 0.016865982485717, 0.184992314547056, 
    0.158968554431872, 0.0129476274228285, 0.132912110415635, 
    0.0191968521890393, -0.0641676508427933, 0.759179972775658, 
    0.262133884769608, -0.0358592699322605, 0.402828462394859, 
    0.294947688342937, -0.0509596342722093, -0.11877777726022, 
    0.168363284933379, 0.0292995616747459, 0.572184516062598, 
    -0.178329509426887, 0.592557803213784, 1.33615129080172, 
    0.184954888470982, -0.111720647258567, 0.321265465613995, 
    0.684602909339066, -0.169533689014324, -0.126237016503011, 
    0.0260468847754967, 0.202305268745212, 0.0730060183890044, 
    0.0171139016774555, 0.0283834784974635, 0.0775863363749812, 
    -0.0403133387415336, 0.018462379679014, 0.314650242247672, 
    0.161152730693409, 0.0742683427660869, 0.178626322766278, 
    0.175505543535231, -0.0737583498725211, 0.374216301210928, 
    0.279943265937957, 0.0628727088652241, -0.015304165809456, 
    0.272203882593383, 0.277217838210292, 0.182331724115204, 
    0.114523884350198, -0.0556017119908367, 0.260645077415127, 
    0.169617991725548, 0.0840816059316777, 0.285229808113944, 
    0.129260170446806, -0.0552068596265209, 0.0339592056752238, 
    -0.158208306224831, -0.00915550381998099, -0.121476571697427, 
    -0.121658639905502, 0.015596269157498, -0.0583704416444879, 
    0.0371611683412471, -0.132376558563389, 0.0301503244495824, 
    0.127690079907054, 0.0515768291141662, 0.0975467052274794, 
    0.303120964060684, 0.161143583583346, 0.0147544427851411, 
    0.532938038784812, 0.144805714157892, -0.263947498721431, 
    0.213031321809861, 0.488278179928046, 0.0763115196231977, 
    0.136320961225684, -0.316640660246373, 0.629177790851608, 
    0.335130125662675, 0.0398162326210001, -0.104544101168122, 
    0.373503359081124, 0.518483575014338, 0.177183536486288, 
    -0.0947477044490608, 0.192032732197242, 0.362753276623617, 
    0.141578430082571, -0.00621177589460763, 0.374358523249468, 
    -0.00694205279421933, -0.237370200846171,
  0.0482862137043773, -0.150353285965098, -0.0490926815975551, 
    -0.103316982033364, -0.0636664946815306, -0.080320766612656, 
    -0.0296249349523611, -0.0847667169215964, 0.00406232230690838, 
    0.0952973821598058, 0.411842012183044, 0.0663697840364501, 
    0.561007977001904, 0.368233379184607, 0.0913791657989151, 
    -0.322495149321451, 0.624491887859337, 0.360377466648346, 
    0.162521706887705, 0.395502900045101, 0.272848717675715, 
    -0.203967684229702, 0.112170523490632, 0.696990743292077, 
    0.287146908176822, 0.116866336814139, 0.428974674026088, 
    0.278932106475262, -0.0535941811087984, 0.472795558113252, 
    0.524875916416225, 0.206227296707859, 0.0922565096120638, 
    0.0708052039288991, 0.0705815704130556, 0.0653429967004802, 
    0.052234370728269, 0.0400237682416491, 0.0487376735144033, 
    0.189998566228126, 0.195346802186995, -0.100276434785633, 
    0.017852786856044, 0.501677934774426, 0.111443915717508, 
    0.143079655635021, 0.252964636848474, -0.263891253698242, 
    0.334887601031593, 0.485228355334501, 0.173796295582321, 
    -0.469733223779484, 0.199318638392919, 0.681555849625055, 
    0.139905792832887, 0.0222316241780548, -0.0701122611918811, 
    -0.325174304136705, 0.577137874955182, 0.440806165457698, 
    0.102600209585969, 0.225185195485741, 0.156632301635692, 
    -0.0153883992004771, -0.0223987783319293, -0.105675665621763, 
    0.113874291724502, 0.158062139575879, 0.0415737672817115, 
    -0.0894065371324132, 0.0526089052660825, 0.0975470869873818, 
    0.0707653512909613, 0.36485068211023, 0.290218418617493, 
    0.0598248107613186, 0.0281452454939141, -0.184944551378052, 
    0.298328979118219, 0.298768647339921, 0.094965360060224, 
    -0.124740016483632, 0.105828150254031, 0.383018588397312, 
    0.063814300047686, 0.0115103397599504, -0.142068007155665, 
    -0.0689953123446292, 0.425762374588798, 0.139376040189516, 
    -0.0624123744050909, 0.0783057527108837, -0.0756482889621244, 
    0.0558895399107099, -0.175120755784772, 0.034346637696768, 
    -0.243424012607735, -0.0693885818479127, -0.202488653732103, 
    -0.200891443316355, 0.0499366794985762, 0.0267706904059558, 
    0.0730665260130001, 0.0793158751268973, 0.0800440166366526, 
    0.0313020951344971, 0.0427783141858692, 0.0771429361918856, 
    0.0783792529723384, 0.0179149965274304, 0.0606886831202483, 
    0.0941565491792638, 0.109048000724398, 0.13442425056122, 
    0.139338082674653, 0.0928529671722085, 0.0906475696561993, 
    0.2628785545717, 0.156361743878576, -0.129667498869817, 
    0.234706424992692, 0.342684460287873, 0.00887135172333686, 
    0.150616737912989, 0.567469867344904, 0.112250329024507, 
    0.0289314018341524, -0.173886343240009, 0.437629654843517, 
    0.309944658834129, 0.0683797377593065, 0.337350176112364, 
    0.400825719800642, 0.121528517760189, 0.752393301997808, 
    0.344113648576748, -0.0916416750233034, 0.459085140308514, 
    0.396383657626792, -0.229951482734208, -0.192171394588393, 
    -0.0448260765042883, -0.262206140860255, -0.0967785626454982, 
    -0.219813225015991, -0.180331680746984, -0.171345069658676, 
    -0.192585914656212, -0.0883940390229938, -0.185853118417476, 
    0.0876293291975937, -0.0523337417874588, 0.0365502998983458, 
    0.0341109275056644, 0.0636124843988063, 0.0261250090579119, 
    0.0723217690237164, -0.0100853784274667, 0.0516921284840103, 
    -0.0555911074165186, -0.00907349164666339, 0.0404856049511702, 
    0.056449118074262, 0.0642693752377909, 0.123437877321968, 
    0.0459087530914955, -0.00576191594375636, -0.00588619977058211, 
    0.214667685774525, 0.0240227282765831, -0.123228747494751, 
    0.729445115941141, 0.537410041251999, -0.340444961709311, 
    0.493932056942749, 0.724546401111673, 0.0736131144829538, 
    -0.200223671020219, -0.021324808808275, 0.901560183420932, 
    0.0504787503788587, 0.0286129231034413, 0.0989603358498289, 
    -0.0102975552903802, 0.0512470295610613, -0.253705552923164, 
    0.289004645914826, 0.160057687279036, 0.156612149972894, 
    0.160875407419587, -0.0208805819888931, 0.112482440950294, 
    -0.271993121559341, 0.0557802971178406, -0.387650079369738, 
    -0.176308515746342, -0.0583272777257439, -0.111061695996465, 
    0.0377599411206557, -0.301004703687747, -0.101008760275523, 
    0.114479486528907, 0.0258462848633931, 0.145421304508452, 
    0.220615969519791, 0.135506002397702, 0.145524095648905, 
    0.0156729836635681, -0.0534413784726161, -0.464550049724721, 
    -0.0513170159439907, 0.614419159248617, 0.373738892691654, 
    0.241520350001183, 0.454140512909688, 0.152086587874039, 
    1.00559176988778, 0.378287272042331, 0.0137048570440463, 
    0.0771327421229762, -0.304594591020224, -0.169487818610067, 
    -0.190921005004664, -0.0920203443045133, -0.205458758184021, 
    0.0416204615766303, -0.282972668511564, -0.052221029580526, 
    -0.217195710321798, -0.227437920554936, 0.0197223914530559, 
    0.0812126768168745, 0.0817173149306158, 0.0861967289882901, 
    -0.0375162879563624, 0.0553969539026627, 0.0141779011039396, 
    0.0954341102936986, 0.162249443049858, -0.043787395652976, 
    0.0199347251760692, 0.064472743834531, 0.0786077967909937, 
    0.10015874584609, 0.114664004248435, 0.0873945066481525, 
    0.0773714333983119, 0.19019592739006, 0.151647196164145, 
    -0.154315069748933, 0.205434905722011, 0.367908205601831, 
    0.166169022315712, 0.127981253448267, 0.257807866597861, 
    0.101041659856509, 0.153558479307093, 0.765931439224949, 
    0.235920817008449, -0.0845550605051555, 0.034251050534993, 
    -0.0452168670124624, 0.827640392422266, 0.0468787629317291, 
    -0.0777785866098472, 0.610721322863556, 0.366195601025714, 
    0.899385813545527, 0.480681396521961, -0.061102103092371, 
    -0.0700169356523807, -0.203713990156468, 0.0942177235121752, 
    -0.208526624394304, -0.0341660239439955, -0.204786043371524, 
    -0.11166139988714, -0.312154812381556, 0.00182017168366634, 
    -0.108114611163622, -0.122456937865795, 0.0807135355918913, 
    -0.125863593954735, 0.0112360497245517, -0.121107803389304, 
    -0.0185896099618461, -0.0761076639109935, 0.00472777251974076, 
    -0.107114518783731, 0.0605597705028605, 0.305846336628702, 
    -0.0400006915605255, -0.214434644848477, 0.573035202043968, 
    0.329079172833724, 0.0967263405128051, 0.454480616860553, 
    0.295394417256862, -0.0691433599321099, -0.139595247035875, 
    0.484203429074071, 0.407150713091117, 0.193850754180471, 
    0.126238470713257, 0.103787261661517, 0.117416984847994, 
    0.159309658540071, 0.126934757053132, 0.0615553953962702, 
    -0.010079903134966, -0.126366879286464, -0.0996329052553969, 
    -0.0148080867819638, -0.0994033193521075, -0.00292999813543632, 
    -0.0596317131494523, 0.0166713547394984, -0.0979344401667904, 
    0.00644083351835673, -0.164747149848895, -0.0380194034376515, 
    -0.0614605780272503, -0.0788720134990244, -0.0481878537525873, 
    -0.063527013040348, -0.052255896463723, -0.0233846829590114, 
    -0.105459151254872, -0.0351014092277548, 0.174679340681487, 
    0.185799143984584, -0.0491791151637441, 0.475396655471989, 
    0.240498143013197, 0.0464820103684465, 0.290700499622099, 
    0.48715455223247, 1.13637398154693, 0.594401559803103, 
    -0.0479769119485942, -0.130187106802606, -0.0127601666894494, 
    -0.0023134574901915, -0.0186532845438382, 0.0337221619848758, 
    -0.0602207005666254, 0.0182007520370917, -0.0436953436533195, 
    0.00276226991116316, -0.0243784643833952, 0.0157354456654964, 
    -0.0668529865443018, 0.0369373822783637, -0.0316300002475847, 
    0.0255020636608459, -0.0860411550618425, -0.00395619575370049, 
    0.000485997359283813, 0.0518953595098921, -0.128760337942157,
  0.0406321244090588, 0.080350301947952, 0.0998573153352583, 
    0.132560855284045, 0.153456626642815, 0.118671264223017, 
    0.119687519008379, 0.217718789280355, 0.135629265082321, 
    -0.0392145491636059, 0.0522200111906293, 0.453037595276253, 
    0.189569338520598, -0.130750629168882, 0.171655164100661, 
    0.533428048553067, 0.112086951718022, -0.0947106414839842, 
    0.00243972024117062, 0.560118076605693, 0.130311441301871, 
    -0.203551161529963, -0.0927174533838191, 0.677490824543279, 
    0.316106784414476, 0.0478722192462333, -0.148249718046607, 
    -0.174138725857138, 0.505618910687271, 0.397189148367228, 
    0.204936145741382, 0.199135603243968, -0.0543041464072481, 
    0.114323103031182, 0.399831249516796, -0.146302690114251, 
    -0.199090580494394, 0.0660612541020819, 0.2297725507333, 
    -0.0618369245088721, -0.00183728240422379, -0.209087612764417, 
    0.0921253751282597, -0.124672731899686, 0.0783361324667635, 
    -0.196323986257402, 0.0675841603093229, -0.226155960468283, 
    -0.00574691316872608, -0.240160084905653, -0.0646434559247688, 
    0.00913996608508944, 0.103236926764644, 0.24946512758276, 
    0.151115176030241, -0.100694276551685, 0.0945428103666724, 
    0.429267274148761, 0.170652093218797, 0.258341677988663, 
    -0.25281348068792, 0.45986615974275, 0.564231868271249, 
    0.109800635964447, -0.113057542299534, -0.268810917812149, 
    0.449170696633634, 0.514528187729163, 0.234371578182914, 
    0.172035131448491, 0.491607681175928, 0.270036313361406, 
    0.239119038686961, 0.225776819200852, -0.178361584781524, 
    0.38948781639595, 0.214719370323495, -0.112175217954459, 
    0.134427364638767, 0.446925051958089, 0.108264142161989, 
    0.0437316110665811, 0.0381910369938099, 0.0602600951666879, 
    0.085433625308099, 0.0560850165181851, 0.0182034442625151, 
    0.173227072928811, 0.0350236169270098, 0.057440657559593, 
    -0.232057476782687, 0.225927915943434, 0.414119819531975, 
    0.0974599629124201, -0.0584452512574836, -0.175963446199407, 
    0.349811053148052, 0.350917373174028, 0.21415533483956, 
    0.239726061749211, 0.218128042889281, -0.21081790841481, 
    0.397441971081266, 0.288663581996866, 0.304618002332122, 
    0.437810418690186, 0.0809095547397742, -0.0102785209730517, 
    0.167768750661258, 0.274640420082776, -0.259163271341677, 
    0.387241036978726, -0.21756323172259, 0.190184435618248, 
    -0.475438176529714, -0.0249466319130637, -0.236425502382514, 
    -0.233161060193084, 0.29794682008494, -0.493946471921966, 
    -0.0110813459802829, 0.0390470489548036, 0.156317995710667, 
    0.223572823401314, 0.199316868986333, 0.13045844670244, 
    0.094794026449122, 0.109401661869671, 0.171904684746939, 
    0.197344522289875, 0.12926851691781, 0.0648861939966973, 
    0.0708026551741876, 0.087790225020392, 0.0770057089448913, 
    0.100149823159199, 0.106273733750354, 0.0893552281214428, 
    0.105107921815446, 0.0784740136894751, 0.10795837267093, 
    0.116388826618938, 0.11951654304144, 0.115653312452125, 
    0.0854033465395513, 0.132492221431218, 0.225759311989715, 
    0.126250687327421, 0.149912315574536, -0.299094603655768, 
    0.371545900579704, 0.443556696267527, 0.540794293622856, 
    0.220123565404997, -0.299057038477952, 0.065033664328849, 
    0.549435787424155, 0.158593419077848, 0.919744113583553, 
    0.404408917344827, -0.307636836932914, -0.193891096008192, 
    -0.0524830461861047, 0.579361031832438, -0.0446159477208513, 
    0.294609294196488, 0.767074917462551, 0.183551194557036, 
    0.188530824194506, 0.899445755917245, 0.227236078765706, 
    0.0339503281734563, 0.022205642436118, -0.153262064985787, 
    0.0670114959462949, 0.191060295384132, 0.0244272912120555, 
    0.0585735248871426, 0.135630334244641, -0.259625620070636, 
    4.25614688820339e-05, 0.433842992679819, 0.180034662675097, 
    -0.112673990447565, 0.198206733643428, 0.350408985246672, 
    0.0947796000450087, -0.0676596579510775, 0.0928698172204582, 
    0.488335853769227, 0.21643901342609, -0.00613700083332532, 
    -0.0978580491493803, -0.0276912485401423, -0.0687958644435682, 
    -0.00117077442770699, -0.0447076943719713, -0.00829891767465579, 
    -0.0749889830350023, -0.0558684770325925, -0.00872064296651008, 
    -0.00264319385632773, 0.0496449373947575, -0.0505058462598375, 
    0.0229098757030832, -0.140408939315156, -0.0428626445312413, 
    -0.0263450213663047, -0.0526113536154403, -0.0624582187860219, 
    0.0428097187293703, 0.047264177305114, 0.0604131091655065, 
    0.0787574435368576, 0.0905780649327994, 0.0653170288624351, 
    0.0608286895666921, 0.0907126763821884, 0.077463538785965, 
    0.00626696025488932, 0.123790833879486, 0.181007689145781, 
    0.105447804290698, 0.117688257161492, 0.284334104578047, 
    0.267028467512703, 0.202853246083678, 0.152828960487318, 
    -0.0343934017231491, 0.218628094049909, 0.627430683813604, 
    0.0854019787903636, -0.14238269899442, -0.151365605893878, 
    0.478041991741607, 0.451291337197563, 0.210673756276292, 
    -0.130577635403194, 0.395220817752251, 0.357139575515723, 
    0.1511134809833, 0.103072035074401, -0.15985361580672, 
    -0.00995480873354355, 0.279901986061649, 0.150468371938895, 
    0.0495141322618765, 0.412596931490666, 0.162529324808823, 
    0.0427804238167249, -0.158603218413665, 0.198006534811793, 
    -0.244603271833613, 0.126691689692848, -0.323811838445207, 
    0.0151161026242986, -0.283833436245983, -0.0756595325368294, 
    -0.198071842011718, -0.132405964939186, -0.0239388424854158, 
    0.0794919270644836, 0.0590901269843625, 0.0802850990904024, 
    0.0746244941213287, 0.0573602321068998, -0.0158288819933268, 
    0.036572713522791, 0.0651517260075251, -0.00871861610275569, 
    0.0827969405362734, 0.154130823088932, 0.0893586601955962, 
    0.0648072459294614, 0.235346677557901, 0.261049866302065, 
    0.17371214414913, 0.066399804948717, -0.123308320155262, 
    -0.080819770567376, 0.454929785693141, 0.264404720289235, 
    0.129255326499263, 0.0801397104981142, 0.0314927439626707, 
    0.413426377529209, -0.00851081880642275, 0.232733359001213, 
    0.976425414926258, 0.244988540551732, -0.0463784815628826, 
    -0.0752229214574375, 0.155099415873121, -0.0250374470996861, 
    -0.0689177810399981, 0.0785579003387677, 0.00265560523509787, 
    -0.018211324185359, 0.024993813772333, -0.0733806979018662, 
    -0.0798239975249268, 0.0380130365673167, 0.164682575568393, 
    -0.0932697159731878, 0.265503596999786, -0.339896147313779, 
    0.0672559995090181, -0.169805446760559, 0.0999913886470022, 
    -0.259068605464241, 0.0190706088491103, 0.0421133866115573, 
    0.0659633840542873, 0.126209977390322, 0.147264602179208, 
    0.120793408610842, 0.124544488620539, 0.174986237447915, 
    0.132322616407606, 0.100715779597907, 0.277574001411217, 
    0.191173214935422, -0.0265573890176656, 0.334101105947011, 
    0.560510180701893, 0.223320225491897, 0.0523057854123721, 
    -0.187869515700612, 0.300004626018843, 0.677379176953373, 
    0.125951540504334, -0.0988779521586629, -0.14113594801745, 
    -0.183010740430239, 0.74187938534182, -0.0645298384976583, 
    0.0464939001947412, 0.397679512968527, -0.389549879523054, 
    -0.0844533133922855, -0.260918709788655, -0.0751419350171421, 
    -0.332526443732856, -0.116625765167075, -0.266215924976093, 
    -0.143407678875944, -0.234015960923848, -0.137296384419574, 
    -0.177704536895733, -0.138424284972157, -0.0277239693362993, 
    0.0899404891582382, 0.0368703303640332, 0.0466877688685967, 
    0.0955951636722477, 0.106494731799382, 0.0143047339524657, 
    0.105839520921558, -0.0141501641389749, 0.0172563047405462,
  -0.267419203363924, -0.0792007793034742, -0.0767525212045316, 
    -0.103305989452676, -0.0561162729347799, -0.0842442014077865, 
    -0.0848491839128636, -0.067349993899373, -0.0558670943270251, 
    -0.127177246820565, 0.0319264328984376, 0.0918037777310493, 
    0.111766393128206, 0.120715853094741, 0.117419569935803, 
    0.0874430801236261, 0.109422200800667, 0.21692376428214, 
    0.100888469209824, -0.0544428209322674, 0.152554337225828, 
    -0.141620278350265, 0.404942248808142, 0.602274537014933, 
    0.159244008780134, 0.0167562316937893, 0.0187899099452515, 
    -0.327412464636324, 0.695225332077219, 0.298197091982931, 
    -0.128064323610821, 0.319265536564081, 0.617924357618406, 
    0.192665378791354, 0.0461193393019424, 0.655066272764364, 
    0.131369857779652, 0.0219209287529898, 1.06628795031589, 
    0.252449821924626, -0.0237801264336419, -0.0290414258066609, 
    0.0465812564747837, 0.0474461731872308, 0.050801719076276, 
    0.0244717576432454, 0.0095055717859974, 0.0947786157279871, 
    0.173285668730615, -0.114697236217234, 0.401317421968164, 
    0.312139591661574, 0.0819210773931519, -0.216894889819721, 
    -0.0191567341281304, 0.471783640708577, 0.378722821073371, 
    0.137751467873068, -0.105180743552137, 0.117378270137577, 
    0.188903728420745, 0.0553369001700984, 0.648133097891956, 
    0.394415119036411, 0.0822269191487677, 0.0808141551907269, 
    -0.235407550828758, -0.089964995693391, 0.384583851770014, 
    0.306321626408304, 0.129669798205953, 0.26455517843161, 
    0.384599353374216, 0.273284699140331, 0.156309338701239, 
    0.132108724634999, 0.194197047801955, 0.176251857947096, 
    0.101072519775889, -0.120549412256402, 0.362814580360982, 
    0.260167742834358, 0.0628971851989006, -0.0332039849096076, 
    -0.0940162434122399, 0.372153049780332, 0.247629407670414, 
    0.24931038804426, 0.54161761651163, 0.197681387691712, 
    0.0285462284329588, -0.178402098135969, 0.0218803296240017, 
    0.600371769515129, -0.0513735174410006, -0.230753345155691, 
    0.0378969762952585, 0.378734061868264, 0.0054674491634428, 
    -0.014764184092362, -0.389034646059578, -0.120925900664831, 
    -0.294035525503297, -0.17428487902565, -0.280505497848662, 
    -0.145049438737015, -0.263150202515766, -0.142206125239691, 
    -0.190602824296926, -0.167925156928052, 0.00559830736360534, 
    -0.065304252611033, 0.0300097041680097, 0.107906032388532, 
    -0.0101726488997255, 0.108187883532139, -0.0670080224491896, 
    0.00356938281695085, 0.0346217372614636, -0.162036444633936, 
    -0.0190194322042461, -0.0438019309732195, -0.0441068096920395, 
    -0.0478764110885763, -0.0132859337042444, -0.0426023121657986, 
    -0.0460096108153678, -0.0119388851347585, 0.0937790309161089, 
    -0.361312833661127, 0.2594232232041, 0.447395952303032, 
    0.365260428438829, 0.179302300891927, 0.167128303509026, 
    -0.4187212059522, 0.352343531205692, 0.532120344324233, 
    0.329930328930931, 0.0413107817653614, 0.277350159850938, 
    0.240456165563031, 0.0834883606262648, -0.0448392043478265, 
    -0.102779543590097, -0.205892559137979, 0.140899543353143, 
    0.123602517646702, 0.302843862080713, 0.120770896327916, 
    -0.186110157240323, 0.0729037850754356, -0.10687351891774, 
    0.108473086405178, -0.572033947912219, 0.00240795603090917, 
    -0.186575394475583, -0.215692539779721, 0.0466250803273578, 
    -0.412395633445099, -0.0734563814797374, 0.0671552775002686, 
    0.140455921672832, 0.132905814607448, 0.110955990135976, 
    0.180608822585471, 0.290266159107278, 0.283030818125196, 
    0.204782642247174, 0.174255036437666, 0.294953699921911, 
    0.343756946563058, 0.313051657000932, 0.309866234401957, 
    0.361498236789318, 0.376148705054466, 0.360256956950488, 
    0.352081590409113, 0.286565010194809, 0.229060052473574, 
    0.400549564888573, 0.468913800667293, 0.2242084518069, 
    0.0370698739993145, 0.344398369383428, 0.442948045609099, 
    0.201821232352519, 0.0890440418291488, 0.0888514786564156, 
    -0.0405809037242104, 0.26968570944376, 0.788496317236079, 
    0.216601987679444, -0.131059573746386, 0.0127954966873128, 
    0.404192800938366, 0.391213856699789, 0.38032604354954, 
    0.257070697604386, 0.257011814268049, 0.671515019003397, 
    0.23590585763915, -0.0461933424338858, -0.0651408054754434, 
    0.454901064745813, 0.132377243765472, 0.275647582646694, 
    0.534150322312848, -0.0457184505677034, -0.0875316413516795, 
    -0.176004944528061, -0.0781497650746107, -0.0186967887299188, 
    -0.0848666249847529, 0.0791924172539548, -0.145006078962174, 
    -0.00771823562738862, -0.00321210813505472, 0.0437801144925317, 
    -0.170382363494221, -0.136357234695236, 0.353916161005125, 
    0.121483733563031, -0.158328512222668, -0.00533246693341347, 
    0.489637671601915, 0.20199249321603, -0.0463652579901306, 
    0.28059725196044, 0.29194600977701, 0.131879692636458, 1.05882324296757, 
    0.261789882011157, 0.055476334466576, 0.535097258137889, 
    -0.689924807344032, 0.438576819488547, 0.71933424580621, 
    0.253384859059448, -0.12177234513202, 0.487976317132629, 
    0.350849214736395, 0.00513980443977739, -0.197528444025182, 
    -0.0297043087955556, 0.611860404551239, 0.103725626233238, 
    0.0161626313167872, -0.175981014382295, 0.00907293785881734, 
    0.344758788919596, 0.222887246919991, 0.0679602445597923, 
    -0.256066476145618, 0.219356251903341, 0.237552877435829, 
    0.0583862949759974, 0.0320166367881773, 0.264918915779767, 
    -0.0622590440756051, -0.0694107394938875, -0.161106449885233, 
    -0.0553342840691998, 0.0599131779225713, -0.0337432477337449, 
    0.0199242937324737, -0.119921262016388, 0.000485616899346564, 
    -0.0698535944115327, -0.106630639166862, 0.0533953533876783, 
    -0.102280492036836, -0.00236519449734711, -0.072960600168822, 
    -0.0279455806534905, -0.0491375697663349, -0.0346698119120901, 
    -0.026143842382433, 0.00562008903465359, -0.0476895730687713, 
    0.164601384702108, 0.0335180542430049, -0.076722597819, 
    0.0410753466899808, 0.439636719975159, 0.169518688135957, 
    -0.0991506548029499, 0.137610471325209, 0.429654028676863, 
    0.210511507544285, -0.392168287139473, 0.251635396154664, 
    0.44391348741477, 0.0821867141958373, 0.757027717575434, 
    0.712911634909686, 0.122980718529523, -0.26819480330251, 
    0.381594613072702, 0.51432573292792, -0.154455549161713, 
    0.050908265757897, -0.254334411275862, 0.014097056822389, 
    -0.261431391446099, -0.132271244935274, -0.0529133223572652, 
    -0.13074356589461, 0.103465133278379, -0.224784070958473, 
    0.0249178771614644, 0.118859713110417, 0.154645330923022, 
    0.15380406196131, 0.148586459811283, 0.147790569497063, 
    0.160589011437376, 0.169111960206252, 0.183388658875939, 
    0.151582341746998, 0.141372164216141, 0.144717093197754, 
    0.164524826636311, 0.190531341533396, 0.192890659298274, 
    0.179448678798093, 0.19402014455995, 0.22618264160187, 0.217043890542722, 
    0.199357487314944, 0.20480669207993, 0.180323921436439, 
    0.164310640771332, 0.261562851248692, 0.279821995678747, 
    0.147156802600151, 0.118423089230351, 0.383282298092676, 
    0.261914323886963, 0.0594964902804938, 0.231515406866049, 
    0.375794600013436, 0.0542061885387627, 0.17129021034968, 
    0.740413541760288, 0.163469779483552, -0.00270858008611928, 
    -0.101222037929265, -0.10419476130523, 0.527988300693394, 
    0.533033059661453, 0.090885279007352, -0.0213679630448629, 
    0.245292978553294, -0.275689564209137, 0.461804917787415, 
    0.456146376630417, 0.0403482164390276, 0.704005485106427, 
    0.339028122232569,
  0.272300316242991, 0.024444725764248, -0.0338739382083895, 
    -0.0652343544738144, -0.122397820230634, 0.0853324768324336, 
    0.0816330661000683, -0.0747023519386963, -0.215508674788491, 
    0.353851487713544, -0.0628928791270098, 0.242603824025245, 
    -0.193566720943592, 0.180505290455823, -0.149675177010542, 
    0.148879421920798, -0.205729055888931, 0.0270310194415107, 
    -0.373786294997522, -0.174274759878228, -0.0135650068514062, 
    0.092796906889438, -0.0631471973620452, 0.00405817906297128, 
    0.0166453679026623, 0.0403673810588807, 0.00157864410778504, 
    0.0249863100036413, -0.120364837816783, -0.0105965705806884, 
    0.0193446818983791, 0.0691471771221285, 0.0618148039919685, 
    0.0281580942716611, 0.0873119032984411, 0.0703874984020863, 
    0.146605501831915, 0.136828063830026, -0.0469646366233519, 
    -0.129466549219104, 0.321769070136853, 0.186810007791532, 
    0.762525627809611, 0.079305302313788, -0.0848848209777381, 
    0.00986901470371238, 0.1196782138321, 0.292544557582236, 
    1.05245883072057, 0.248782403817809, -0.137527654626869, 
    -0.0596919375002067, 0.0256300820113687, -0.0280491552580794, 
    -0.0363038820324334, 0.130933814232676, 0.0491357016040864, 
    0.273910905699195, 0.238424344243013, -0.000362987261566056, 
    -0.0182727745069257, -0.0288728910071038, -0.473146460971579, 
    -0.139003122693639, -0.153954516697919, -0.443121556809396, 
    0.156670411015549, -0.194601318403378, -0.0372662135154238, 
    -0.387088498790203, -0.144878786647658, 0.037639347465099, 
    0.099738295346703, 0.134739193659396, 0.139693507400189, 
    -0.00391456596353673, 0.0370444017549748, 0.051544956029294, 
    0.0620417410610253, 0.0646497515520748, 0.0524512236674868, 
    0.082294898068353, 0.0358643545601071, 0.0564754151949841, 
    0.0424151230174829, 0.0376763051849227, 0.0589637740057234, 
    0.0510507929350074, 0.0597018254420005, -0.0211921385660144, 
    0.245979666218732, 0.168114878630232, 0.0355026699827823, 
    -0.0340316617104004, 0.280990511042839, 0.308609172252261, 
    0.243773578110052, 0.225292720118757, 0.138514284043104, 
    -0.410132337865198, 0.190125525684615, 0.569010420450425, 
    0.481192464010939, 0.322101486786848, -0.0645938355166329, 
    0.726947687111524, 0.318848381134246, 0.0655513835330669, 
    0.1464541515011, 0.643642095819709, 0.109535794727613, 
    -0.0101395554827305, 0.607561748255136, 0.399308903124551, 
    0.070010886349775, -0.124903354223576, -0.0183937012968404, 
    0.272309412401936, 0.235799231273743, 0.294716935244063, 
    0.263001272313096, 0.0700257887214284, 0.0157371985112271, 
    -0.0178182229030559, 0.188252503071963, 0.0408945705141878, 
    -0.093151650442605, 0.0372250203163275, 0.179469599020872, 
    0.0745141339348, 0.0691404134849148, 0.205775891604361, 
    0.199662073801369, -0.00919663526148767, -0.0221287579133468, 
    0.455160088678922, 0.196582120452044, -0.0173416014696798, 
    0.287889009372819, 0.337560365797168, 0.142741396492734, 
    0.0929523158250082, 0.0808354229419894, 0.0884943819566344, 
    0.0788050849210609, 0.0863480636892823, 0.0599431508760954, 
    0.0673984845750583, 0.0780453866607196, -0.000721233586928244, 
    0.297115507624347, 0.206099336878441, 0.062191272473457, 
    0.0353689695421665, 0.171981249589158, 0.582381188730083, 
    0.246520001858728, -0.0374602039711786, 0.0259330966248943, 
    0.375092722313192, 0.353939127154616, 0.20350353156347, 
    -0.0233625025614749, 0.438064949479912, 0.858050282347405, 
    -0.187887482240366, -0.19541761149704, -0.00214961905495384, 
    0.741244304416417, -0.0543602555490277, -0.0540001514997437, 
    -0.249323671858574, 0.0526288424295563, -0.264991575571877, 
    -0.0254966963491561, -0.22706106129178, -0.0372501505670182, 
    -0.181494552091462, -0.136991014203478, -0.061415074314932, 
    -0.100864173378466, -0.0110930613975828, -0.177680475886632, 
    -0.138669623552092, 0.168839559699928, -0.119209182170345, 
    0.0850118137643937, -0.0256132311710934, 0.0388365295354704, 
    -0.195489325419426, -0.00761265697468823, 0.0897861161949027, 
    -0.00382868815518217, 0.0728112132012466, 0.259013200671452, 
    0.10417130910268, 0.129543251244864, 0.260092030101413, 
    -0.263604394286385, 0.368386124735704, 0.316352387107551, 
    -0.00469618071270643, -0.310675174645574, 0.133333615837707, 
    0.758682769337018, 0.369666701896061, -0.0988561629636229, 
    0.307181006632779, 0.522256267522344, 0.37309042773022, 
    0.286531260345824, 0.212530138662465, -0.070252591961114, 
    0.808405731725281, 0.26749764448861, 0.0218146403719868, 
    -0.173389283608414, -0.132716823429435, 0.638424284063034, 
    0.289585656229624, -0.00914622572329144, 0.124919237668645, 
    0.0965541644983691, 0.220053254343813, 0.0388805039469121, 
    -0.207777048772336, -0.0956873296483077, -0.152536815827326, 
    0.0855297013317552, 0.0421091304492897, -0.291310390750239, 
    -0.016339695971742, -0.174609302993189, -0.0303277432584259, 
    -0.165592663465175, 0.0717157003233379, -0.141608405112422, 
    0.0713236938664157, -0.278738601534797, -0.0880063212201213, 
    -0.00383690692130792, -0.0333805647663333, 0.0642195285459172, 
    -0.0251627135612413, 0.0516522862440974, 0.0135861304289246, 
    0.0460442007409686, 0.0218429799533698, 0.0469724612207236, 
    -0.0585476750729546, 0.0399733192917044, 0.0313991990613421, 
    0.065936486808201, 0.102948211388819, 0.0711478700136528, 
    -0.0123457017230166, 0.23058359402557, 0.074854873480289, 
    -0.161470911542483, -0.150989695246343, 0.510091222003126, 
    0.0721833645231551, 0.338972652074847, 0.696876871945373, 
    0.140542438232786, 0.000916400778725943, 0.370237443331271, 
    0.493078833340463, -0.110240329881074, 0.736646176141313, 
    0.346786112861212, 0.0102446003646539, -0.0383233955799255, 
    0.0812210986427876, 0.172233614852467, -0.0306461368073927, 
    -0.0387225155185189, 0.0331917604636572, 0.150939505533135, 
    -0.0308849274886812, -0.0505890874760951, -0.13187484843332, 
    0.0251196975222925, -0.0418192731019484, 0.0529526525290602, 
    -0.104164291947319, 0.0303678729922472, -0.192166875371361, 
    -0.0747130212585897, -0.0349934477530411, -0.0460047631918209, 
    -0.0217845967559091, 0.272423155873579, 0.106341501788345, 
    0.0211012450533173, -0.113346927992479, 0.0331746565400421, 
    0.239278887658415, 0.122033770476322, 0.369481544745686, 
    0.482183365948314, -0.112105654989911, 0.683785585958508, 
    0.573630067935827, -0.0492207334735187, 0.0970801968784674, 
    -0.539621692564668, 0.535008414093505, 0.761557903309956, 
    0.0375002766612035, -0.129635392326812, -0.173477592389256, 
    0.157520667558241, -0.0186526910317285, 0.113788496779475, 
    -0.222800146626562, 0.0578431399657617, -0.154881203581625, 
    -0.0142543704488399, -0.119340988020699, 0.0125087284832149, 
    0.0915701895140745, 0.204087944569276, 0.187309311613573, 
    0.240233338279355, 0.394949396356328, 0.266295115940492, 
    0.0649128849249437, 0.211243074041385, 0.457124772805423, 
    0.301451414153434, 0.200662078603109, 0.174678841974204, 
    0.146505434132453, 0.150492722159434, 0.127094774009105, 
    0.118046709349355, 0.167119343030281, 0.168045800592395, 
    0.093628472383308, 0.101467178049162, 0.225636681655513, 
    0.170688377967327, 0.0620568719372754, 0.145206063987778, 
    0.231543680478299, 0.284165135863791, 0.325931541463879, 
    0.0840215975566453, -0.0714352475124112, -0.291948378777676, 
    0.025293112529425, 0.625514617617051, 0.445430265844282, 
    0.183385088197027, -0.108954485060579, 0.343772871257816, 
    0.039775305997559, 0.124499959628064, 0.927482889401712,
  -0.0768579142214691, 0.0639619556004039, 0.291259030961084, 
    0.398807474240364, 0.355496371349224, 0.192730627679337, 
    0.103351088229776, 0.34010889834174, 0.252779900407559, 
    0.0321925441382608, -0.169170803798654, -0.0526062814310379, 
    0.414200230098822, 0.347388241370977, 0.0749544665344061, 
    -0.129196470065142, -0.0716122183616495, 0.292407343788085, 
    0.188758306143068, 0.377832700868598, 0.410494167965267, 
    0.149212015402496, 0.646921549454171, 0.384650071958314, 
    0.0173738143509756, 0.367551453590702, 0.549102198954637, 
    0.0581712825319838, -0.22972793721212, 0.64630625235479, 
    0.530533748343557, 0.179836239034354, -0.0219321763387808, 
    0.375688760349637, 0.352709744540053, 0.182984789356935, 
    0.115751037374183, 0.108046885875917, -0.130627580354392, 
    0.143340411180407, 0.273821702201341, 0.253680254024938, 
    0.528729780012239, 0.325681474259386, -0.0244808933490173, 
    0.431877749745375, 0.425850469286081, 0.211323829779693, 
    0.295753250537426, 0.261790545079686, 0.03567898224466, 0.53976911327069, 
    0.362541968610104, 0.0355254653125339, 0.186440227216444, 
    0.450521617761312, 0.119868187253267, 0.0330496895049194, 
    0.510235962489985, 0.207946710342547, 0.0324866400891274, 
    0.0251684235123873, 0.0482280067784853, 0.0448286629581598, 
    0.048949926260495, 0.030761551727011, 0.0317447250946475, 
    0.0638473866201514, 0.00398704278239752, 0.133704476863442, 
    0.32079603746589, -0.013092301197646, -0.0384590802869127, 
    0.409171240706016, 0.326869400254505, 0.175807015546594, 
    0.269649026589685, 0.275388301992076, -0.118726185322795, 
    -0.176617057205875, 0.517729354233922, 0.687656106018009, 
    0.0722900017353293, -0.18724087672582, 0.0595297207645494, 
    -0.0186210518646572, -0.179261416034129, 0.570494139409254, 
    0.841541994365283, 0.0220426200980094, -0.325115426447801, 
    -0.0246217546924717, -0.231393600806842, 0.122929124337409, 
    -0.272851934902387, -0.0684381186678463, -0.212305523476712, 
    -0.170409475008767, -0.220400617867087, -0.130350020897874, 
    -0.129259092238016, -0.0504081209159106, -0.0940742698612431, 
    -0.0404748898113184, -0.0325650034647634, -0.0496967040118534, 
    0.113007604240278, -0.0488055333598179, 0.113291366847344, 
    -0.0496590004414948, 0.0373408872350177, -0.0870721052971973, 
    -0.0123797637334306, -0.0575047178752953, -0.0216819320213455, 
    -0.0453241203483603, -0.0512439368603204, 0.0557340615902145, 
    0.0174064683234101, -0.078594117483009, -0.19987523142282, 
    0.111939445601554, 0.379776169463072, 0.0905994386917465, 
    0.0306898054149161, -0.134621221785732, 0.288865565862694, 
    0.281366407149459, 0.175445179137279, -0.00652535111500099, 
    0.504536827201419, 0.215918291303776, 0.135095788323412, 
    0.876742481573593, 0.309623590971873, 0.0879449415405759, 
    -0.0818639730728983, 0.51348354998091, 0.358372223600681, 
    0.0810491049628615, 0.168747493650509, 0.508234907723972, 
    0.393956028291651, 0.240824995684394, 0.166002931401456, 
    0.104355071899972, 0.101630459518007, 0.158421520265075, 
    0.116079402846171, 0.20082262845687, 0.210008810504478, 
    -0.0278818008692007, -0.0223422699248641, 0.444821855519643, 
    0.199073205930277, 0.131307089440833, 0.190794617792842, 
    -0.241063214958365, 0.490631534325091, 0.197314578167121, 
    -0.202587466585505, 0.0774806999712896, 0.620289334447173, 
    0.169637630278475, -0.0996842040755915, 0.216624814955956, 
    0.593174938193895, 0.0461150367453559, 0.120786027656311, 
    0.0452558474180895, -0.447394036896272, -0.164758668784859, 
    0.0164205481276432, -0.228778027154762, 0.102883742688505, 
    -0.155484157161604, 0.039589196044643, -0.0735605365779384, 
    0.088331695242281, -0.286989253543521, 0.0246241054077012, 
    0.0773581830819038, 0.0984440047196133, 0.14120365283242, 
    0.138826688952501, 0.110681006871191, 0.129562654321021, 
    0.0524988791774984, 0.0672975183798395, 0.050102899408323, 
    0.132464142617347, 0.138747361038059, 0.173244982142714, 
    0.18592091381251, 0.17162863412302, 0.103055367210965, 0.2415588353039, 
    0.353282621923213, 0.126188164027067, -0.0639808693095671, 
    0.138207384185384, 0.721630874121667, 0.177643634016064, 
    -0.149810502670413, -0.321336369959873, 0.581877523580811, 
    0.453790734673279, 0.290652852251779, 0.402734805671215, 
    0.146810486426439, -0.105238136683332, 0.717974424434877, 
    0.561749287662633, 0.170426525364744, -0.175701108203777, 
    0.416702292803682, 0.281753170826121, 0.0991884193628963, 
    0.523853800576191, 0.218800680479524, -0.0604320702042692, 
    0.0186336500669862, -0.114856791220132, 0.0679939709225936, 
    0.103758308916226, 0.0195091252423871, -0.0206372479577371, 
    -0.00520461613356578, -0.149134403647088, -0.0496018802923128, 
    0.236026177766531, 0.119248191049034, 0.0268124608711656, 
    -0.0898556106827831, 0.162433987213434, 0.328895619054001, 
    0.131069463871905, -0.0741068591442907, 0.139166439647572, 
    0.250800452908711, -0.0300439827741913, -0.025646017976786, 
    -0.101202067446759, -0.0185841738247087, -0.316449425062625, 
    -0.0889098836442225, 0.00266870148065, -0.160417805025395, 
    0.0739575745291619, -0.161222448579006, -0.00591811348929409, 
    0.0466463912884339, 0.0985912786145132, 0.116726041859821, 
    0.107272366512681, 0.109537480275444, 0.0869048457892877, 
    0.102457364885081, 0.103803308724882, -0.0405513854371712, 
    0.163874700353266, 0.328016821827408, 0.199758884018859, 
    0.0447511788398564, 0.220483302621988, 0.461408938983163, 
    0.212331566207546, -0.0215433658804452, 0.473027095104372, 
    0.478259554413315, 0.0909992269374079, -0.365658682019068, 
    0.0246323982895055, 0.937455369095423, -0.0476421851863302, 
    -0.00320023661011383, -0.113360266198759, -0.390205759157467, 
    0.392841811000433, 0.596979489043125, 0.114148530350767, 
    0.01828903691813, -0.0378950418741563, 0.000361476954209544, 
    0.0666843375962814, 0.0793477160317307, 0.176474457143818, 
    -0.24107549402385, -0.213228989530964, 0.119466073036723, 
    -0.20039221792262, -0.11256674459905, -0.313561984017608, 
    -0.328263110310437, 0.182941689037665, -0.151636298809185, 
    0.095466029284751, -0.0598443510032399, 0.0116635035694267, 
    -0.32477127364078, -0.0689481927687549, -0.00728428364211045, 
    0.00878079478845169, -0.0139439013744731, -0.0639374296125389, 
    0.108101614114134, 0.0344724094881271, -0.0432472470155979, 
    0.120229177738091, 0.0504536540130813, -0.167306683218213, 
    -0.0972109004507426, 0.755279126117855, 0.363190066800699, 
    0.244868655265153, -0.375199322649481, -0.122603882648611, 
    0.587539328203919, 0.373122793158951, 0.150027405787033, 
    0.0176383203455414, 0.375713050390606, 0.173073658528803, 
    0.057913612664708, 0.189039819473185, 0.145575857250896, 
    0.0419234092673924, 0.303179401127171, 0.182538713148114, 
    0.0122821558811067, -0.059501515797537, 0.00416324993270381, 
    -0.107767881219151, -0.0249802244116904, -0.062965152246191, 
    -0.0731660320459322, -0.0219357503654639, 0.0398143028223021, 
    0.108098654321478, -0.124121920012419, -0.0198942870649236, 
    0.0499452103399438, 0.535045785496817, 0.104331785854101, 
    -0.130202708970017, 0.0513570578156126, 0.429461903168412, 
    -0.00410204159592933, -0.121338062814238, 0.0172889515020042, 
    0.487043906614158, 0.269588752785947, 0.144117744758048, 
    0.78414963100586, -0.00938329520098293, -0.698508451876733, 
    -0.212896076142956, 0.990047897671883, 0.504241720774753, 0.16069655189465,
  0.152965720286829, 0.00565584434530267, 0.115174864820663, 
    0.185432070943556, 0.0580338002415606, 0.0731253448939308, 
    -0.0153015151642017, 0.215594011848724, 0.138774733100924, 
    0.227839652394118, -0.28907462614961, 0.240156477867934, 
    0.205106367702742, 0.181660093067663, 0.989825766815692, 
    0.602453713418625, 0.207758318240604, 0.168975113013985, 
    0.933184861333209, 0.0328159158407683, -0.126398527778781, 
    -0.132531895503419, -0.15646525511882, 0.180411769739147, 
    0.0623253229525379, -0.0583926446795184, 0.212007054707768, 
    0.032633052992577, -0.0821945148783968, 0.0682030337231295, 
    -0.218664371611415, 0.0395897719714021, -0.124866180982193, 
    0.0456991070825785, -0.0972705490465424, 0.0668132100112554, 
    -0.291741368335659, -0.0347018875409718, -0.185515856433189, 
    -0.200502721568095, 0.00792658035882773, 0.0846149503187957, 
    0.0895801736055289, 0.0749840893544315, 0.100901743815214, 
    0.0999868010470458, 0.155711998199795, 0.145066264557316, 
    0.0695165575004872, -0.0169912303920677, -0.0367848115015739, 
    -0.181500513616601, 0.0253479964480145, -0.124717598001098, 
    -0.0368892130174802, -0.0143183309482285, 0.0329172124342191, 
    -0.11297670703589, 0.0409003068644598, -0.254892958499698, 
    -0.0607004772254055, 0.00589420120964544, 0.0367840860776477, 
    0.0213529460311921, -0.0155448684937222, 0.0204820494812759, 
    0.0406206310950229, 0.115860965480962, 0.0158343584561021, 
    0.0512326306497273, -0.192688421360307, 0.379119544349021, 
    0.255590446182956, 0.0322660432994293, -0.273823960046508, 
    0.474823240223398, 0.536480807938272, 0.150558007451751, 
    0.172985306539961, -0.224737285455892, 0.657162371223525, 
    0.207799619732002, 0.0495815434498734, -0.0570746556088602, 
    -0.0475953328894955, 0.705266097512281, 0.435174879300537, 
    -0.267179839797377, 0.243662756668844, 1.14061795803687, 
    -0.0250793243090085, -0.0775419106339033, -0.0341654131476278, 
    0.0226060085360856, 0.170962150004994, -0.0977227127460117, 
    0.122354549272674, -0.34312477293376, 0.121784797935488, 
    -0.0859665230477673, -0.211091562020099, 0.0271328129989446, 
    -0.222456391469955, -0.112024025050508, -0.0796311020135851, 
    -0.146683388572955, -0.0240172124970047, -0.112362386928458, 
    -0.0276874227023184, -0.0745934986427942, -0.19158247958712, 
    0.22888361263254, 0.161605052781956, -0.0553060046416626, 
    0.030381454929769, 0.308155123627678, 0.238371625624471, 
    0.192847023872245, 0.0431167151224576, -0.157951627717147, 
    0.00363410302701801, -0.288654617327971, 0.549960946361025, 
    0.430731177347925, 0.334019121163792, 0.802890211423512, 
    0.281455542612373, -0.0542424216812915, 0.50900098745963, 
    0.296528067169652, -0.25524745777516, -0.121788175753396, 
    -0.0187577662765159, -0.225441916499781, -0.0136544493493345, 
    -0.0630544149637736, -0.236689694200407, -0.121719431092381, 
    -0.0474033958433754, -0.0760036970159215, 0.0254073978273262, 
    -0.112917877632187, 0.0826305499363468, -0.199723134612691, 
    -0.0393679266258405, -0.0776724316187131, 0.0127905985755196, 
    -0.0595425867710151, 0.0257650686921082, -0.261645465031489, 
    -0.0241683995720862, 0.0312670079855627, 0.0877019322079352, 
    0.0668233524548602, 0.0667759232491813, 0.0358913947182553, 
    0.0292899671594113, 0.0771822743877113, 0.0652854048996161, 
    0.0177170001437596, 0.073066837640798, 0.0513243651648987, 
    0.044037317724676, 0.0462434281561491, 0.130973465125174, 
    0.0687698658096758, -0.0873177028546518, -0.0523355159033502, 
    0.216341003997669, 0.230725281866391, 0.47858351320149, 
    -0.138519782640336, 0.573382256903683, 0.513723989876492, 
    0.0743333475854277, -0.305955571148817, -0.00149477848598906, 
    0.564517049932416, 0.680683067382681, 0.273457193954571, 
    -0.121548080281066, 0.0582243772702383, 0.762413507053919, 
    -0.0284318484481056, -0.190645667390567, 0.162667124324664, 
    0.408298586976652, -0.0640277431782961, 0.538929154144127, 
    0.560511110288409, 0.055367626597797, 0.0191457266486552, 
    0.0218723670088565, 0.0199606040456929, 0.0257129859432092, 
    0.0268311423195805, 0.00976344998362995, 0.0873706915575937, 
    0.0949438766903669, -0.21786469058164, 0.339784608300089, 
    0.33413339520826, -0.162740007816196, 0.344108985052682, 
    0.53353128179407, 0.0716309871370435, -0.0306093236944364, 
    -0.00118038453251418, -0.258558955977995, 0.633420437583663, 
    0.294555668478131, -0.0687309233512534, 0.151975027387587, 
    0.609357617955891, 0.382874141093792, -0.0871538078560134, 
    -0.146563018201579, -0.400809424815798, 0.131568474048865, 
    0.416767941569326, -0.116935439736669, -0.0877975860635083, 
    -0.398493579726661, 0.00532194503710221, -0.168058937653592, 
    -0.243645742178881, 0.0246527379036682, -0.154300051834322, 
    -0.0731250034751746, -0.143230491920157, -0.203459824678773, 
    0.0576192452771561, 0.460894919280033, 0.167647628623724, 
    -0.283788184698509, 0.162590594986512, 0.53553490506799, 
    0.153368259296899, 0.0331119663839708, -0.0851967134225265, 
    0.0311343052547135, 0.344879780790196, 0.365136243498396, 
    0.339949104894028, 0.411060338309115, 0.328557538329672, 
    0.138545327588855, 0.109156344542987, 0.486475310062924, 
    0.272802158813477, -0.0106047336047872, -0.0110974342980739, 
    -0.0037466638882878, -0.0170637939077872, -0.0111298946291923, 
    -0.0220267813258218, -0.0160689731964332, -0.0191457355296012, 
    -0.0120120264022705, -0.00854270183344212, 0.0229953899421616, 
    0.0118225390880958, 0.042173324011641, 0.010719677696523, 
    0.0273658860853688, 0.0272722342942611, -0.0423512572563157, 
    0.0382084705892359, 0.0570663086283764, 0.0878119057837864, 
    0.126405143442013, -0.0146635206781909, -0.113481948062647, 
    0.321006270143511, 0.46573297368766, 0.23725162455983, 0.100384812192905, 
    0.0717276019973174, 0.127180121089991, 0.0102990406829442, 
    0.386255681075528, 0.374307266225546, 0.0798772093177022, 
    0.895174474631102, 0.477850228436457, -0.0544394106836086, 
    -0.0224727758261515, -0.0240427192780613, 0.505907803312701, 
    0.114087365252037, -0.0302894778581587, -0.0163527896866442, 
    0.0556380439597614, 0.0256743387933902, 0.0715024423443872, 
    0.0117154755035097, -0.0674025845161733, 0.140473267905428, 
    0.0579954685290937, -0.083152777684867, -0.193266575328892, 
    -0.127741492743809, 0.385657334019557, 0.491743493268936, 
    0.198496030805568, -0.139800161888052, 0.0654003131490318, 
    0.534159953535425, 0.437466874444212, 0.129027260938698, 
    0.222887308331436, -0.295118838485791, 0.905953378152895, 
    0.158445744090638, -0.0426240607859027, -0.124309323610872, 
    -0.144150446014798, 0.954117781777532, 0.401923263886285, 
    -0.0242144483454872, 0.236123027670865, 0.556932545810696, 
    -0.0943210551007995, -0.218013132180676, 0.248269180996247, 
    0.179122576864903, 0.0105496319338571, 0.132830320471264, 
    0.0293410115140106, 0.351265831940237, 0.150774184091753, 
    0.0151130898627985, -0.192383004903199, -0.0219826283185837, 
    0.49645421112504, -0.0848132845181978, 0.0631658622488477, 
    -0.079526949363755, 0.388190349994554, 0.11242304510479, 
    0.0304333827965127, 0.0264180698806566, 0.117950205178867, 
    -0.0584886425107051, 0.0948771050154531, 0.0443701349433357, 
    0.040578056368191, 0.346124481693933, 0.0853850283836548, 
    -0.0339707972160438, -0.14589471537631, 0.0215635686138146, 
    -0.133437191175758, -0.0457406893923027, -0.252302872656967, 
    -0.119323467993159, 0.0644894870601065, -0.163950963941488, 
    0.0976427577074008, -0.0225179378842578,
  -0.160193929956157, -0.0524425784415767, -0.0559393130690948, 
    -0.054726115787504, -0.0245834367525215, -0.0577842272997758, 
    -0.0347105017595376, -0.0378646399916995, -0.0606576450128201, 
    -0.0686776237880878, 0.0364903904938668, -0.0106942685369346, 
    0.0562623734962111, 0.00684542487720864, 0.0452161782455717, 
    -0.0299098527146554, 0.029571711729338, -0.00186170106815212, 
    0.0277940890372033, -0.0296124603771197, 0.0213450248871127, 
    0.0403430837002724, 0.0565581579562327, 0.0662091724716562, 
    0.172089034185074, 0.168491429006251, -0.285772889364414, 
    0.276300328948108, 0.40992980662159, -0.270336937096662, 
    0.244678449198172, 0.612698877074138, 0.059940906389738, 
    -0.0246456013748322, 0.819568696065134, 0.590420860209182, 
    0.248396006354462, 0.574109766185544, 1.00773311795847, 
    0.0487485227405421, -0.0900155635730255, -0.0520665982754829, 
    0.188391250595197, 0.0892783227455322, 0.0333329307198938, 
    0.00981978693200437, 0.0883626061065279, 0.0833609542055291, 
    0.02202692578554, 0.00815084456770424, -0.0360749531442723, 
    -0.0053144942002589, -0.0242822348668106, -0.00876540512697309, 
    -0.021145528377602, -0.0143543316297092, -0.00297309811078457, 
    -0.0135774348079293, 0.00514435664024354, 0.000835136684685434, 
    0.0856580741211378, -0.0527160614166165, 0.255266289435821, 
    0.280711262928985, 0.0963752544933836, -0.0404285693738269, 
    -0.0127880008383716, 0.322959597679546, 0.280773472458582, 
    0.146675414550146, 0.191947073111392, 0.315906673090942, 
    0.191260380575586, -0.122537163322682, 0.396331733446712, 
    0.587635638696348, 0.180007634634073, -0.141382586637728, 
    0.489456308737114, 0.5406210289249, 0.06822097435483, -0.226203725994608, 
    0.0696638500396832, 0.532647806865789, 0.145719612401721, 
    0.0489716747623501, -0.159546335999109, 0.180089852822562, 
    0.341834671815529, 0.334752541898019, 0.345530505661289, 
    0.170245963740753, 0.0587291780305342, -0.374553835468997, 
    0.259005459356988, 0.410412192331945, 0.196909867462711, 
    0.0569063440263386, 0.498613799127718, 0.165568125813801, 
    -0.0442223524333699, -0.0736410456228317, 0.0604724186399906, 
    -0.114722309907901, -0.0282259505256097, -0.195901181528418, 
    0.0321363107452086, 0.0176690584416846, -0.0759057275739557, 
    0.119327979399693, -0.286402991329944, 0.0658124970626604, 
    -0.155326496200652, 0.0520938034943731, -0.080015192854672, 
    0.0785046590113649, -0.259555092626745, -0.0446048790336563, 
    -0.181072460206825, -0.192601102190868, 0.00905214229392917, 
    0.056651865261255, 0.0935250618076438, 0.132454483419428, 
    0.13265218841875, 0.125341807489908, 0.164773575820211, 0.19473634950859, 
    0.13443107823078, 0.0635819435044307, 0.139596567480727, 
    0.244564321027345, 0.212652144098537, 0.130846002672442, 
    0.277691570191887, 0.367902677800609, 0.180525877033259, 
    0.110549843267847, 0.460063963929011, 0.309210384274129, 
    0.0778986743166891, -0.01795600848521, 0.482394181897005, 
    0.412016413302739, 0.190587743900327, -0.1874574436275, 
    0.301341657313351, 0.310502583085792, 0.200781873572646, 
    0.525867086092385, 0.287494138009071, 0.0483317635985718, 
    0.0162417818734947, 0.0680868945436506, 0.501284482377873, 
    0.0360414461239399, 0.00374100981866969, 0.338721646072841, 
    0.126737065347036, 0.10260108676271, -0.165304024169852, 
    0.0754993764172696, -0.318676648178532, -0.0543728894402602, 
    -0.171470715528311, -0.196183762146729, 0.0539881246818443, 
    -0.13896660823421, 0.112823590892366, -0.194182170017488, 
    0.0564186401128339, 0.0714920180650293, 0.0853942189179514, 
    0.110978745989261, 0.11250517879096, 0.0667425827426885, 
    0.0775660772028941, 0.112083691786265, 0.102186155642421, 
    0.0402448465251543, 0.101795091178815, 0.14745983337847, 
    0.124377381661316, 0.128047779649332, 0.221133100504235, 
    0.241259434228653, 0.178789664336609, 0.10002594595448, 
    0.0241759203330385, 0.371241449851826, 0.378932748255829, 
    0.0883992428410929, -0.166574029574013, 0.0490948560846394, 
    0.46073518847804, 0.41909407108036, 0.215540302985981, 
    -0.0115226817323875, 0.582502126270646, 0.344196778394746, 
    0.0976050127309725, -0.144784069871689, 0.154433870044299, 
    0.616917472529323, 0.237485834475987, -0.131471899986205, 
    -0.023042213557398, 0.464027173231748, 0.418724588557884, 
    -0.055671697489599, -0.297786728520693, -0.231126682504738, 
    -0.0976484979432596, -0.187195073301982, 0.0311380108482155, 
    -0.197936305137021, 0.106130091459039, -0.291848487386662, 
    0.0439853109420152, -0.161815786185381, 0.129424838139353, 
    -0.0922205387448175, 0.117013237033534, -0.104932768788746, 
    0.0657724950120919, -0.123562823601563, 0.0536648720946891, 
    -0.0652345527407145, 0.0720567734278545, -0.235916451531462, 
    -0.0148889582184286, -0.0120414209439065, 0.0157025811337818, 
    0.0532767568635206, 0.033622235203004, -0.0300306652971477, 
    0.0716524279045895, 0.0798269886452964, -0.0245476792363451, 
    -0.265705665251985, -0.0016499614170651, 0.476858330589861, 
    0.0379373257198049, 0.0460601719672807, 0.616686876186302, 
    0.648265564098119, 0.143589455982872, -0.115622608063346, 
    -0.107508186706751, 0.0559695223262918, 0.622442457600148, 
    0.324026224575292, -0.112027600835329, 0.103561288415051, 
    0.875961834731157, 0.110890795022239, -0.0395248144912668, 
    0.185258299552065, 0.64779251846527, -0.132214463736248, 
    -0.166152203111039, -0.193548270102441, -0.110367135040685, 
    -0.0565345050797449, -0.160988897115078, -0.0395545489728816, 
    -0.235456821189053, -0.0333729088520943, -0.1462111925457, 
    -0.0984196791505549, -0.0538811482411677, 0.146615424176184, 
    -0.0491091303430724, 0.106047138094947, -0.112584145061969, 
    0.0503130370321004, -0.0713056799917174, 0.049250123832651, 
    -0.016078049004446, 0.0594551988639725, -0.104087683986915, 
    0.00353121322598692, -0.0439775816972379, 0.0279193367241663, 
    -0.149569418087128, 0.0245241508261383, -0.0723613095254279, 
    -0.0116122351437128, 0.0857162489648889, -0.149805806165684, 
    0.050217470051973, 0.015333567081524, 0.0394698385355623, 
    0.110118115035477, 0.071232201885341, -0.00339161990626581, 
    0.118971424313926, 0.122202524944941, 0.0360695866361891, 
    0.174274000539652, 0.146872585514836, -0.293522428150331, 
    -0.138407402379748, 0.274417063854819, 0.549241115050753, 
    0.472264376329553, 0.0443213015144639, 0.0811596203388266, 
    0.994064644663506, 0.438371213283758, 0.0759797742856791, 
    0.0929626507876269, -0.000115358036959584, 0.118959526083989, 
    0.026434834537954, -0.0209450649662856, -0.00294029992270214, 
    0.0202498664093085, 0.170440357211459, 0.0997909026624886, 
    -0.0640325359359657, 0.0335697444613748, -0.130669697880227, 
    -0.0316985747975987, -0.0337201388387788, 0.0304682836099934, 
    -0.224142427698879, 0.0186562557367265, -0.283914963553584, 
    -0.192862762405242, 0.0184295646604098, 0.0244505529803115, 
    0.112285567683351, 0.160921084598213, 0.130504330688682, 
    0.096739789518812, 0.0885055771067612, 0.151078295275422, 
    0.146137032777731, 0.0861830212921372, 0.16393027600035, 
    0.235724678014963, 0.187837614503721, 0.133286395372035, 
    0.239969372346916, 0.286990901539201, 0.303284024652106, 
    0.208340297110701, -0.113017679802852, 0.225434087937501, 
    0.488295260559364, 0.0733907735523596, 0.491659966250823, 
    0.635261407837708, 0.101270060141933, 0.278772050306696, 
    0.762431033172846, 0.0368875432152717, 1.02798671642425, 0.659833599057079,
  0.0423958470874636, 0.128399674075654, 0.149676112675235, 
    0.150849739574431, 0.145900903687705, 0.132084986549516, 
    0.153249979369799, 0.198130849948134, 0.17647767071203, 
    0.122315754874426, 0.135301059297058, 0.134859763326084, 
    0.177405315649085, 0.244360611552917, 0.171055363631669, 
    0.0822128541584932, 0.329993218660615, 0.220298859503483, 
    -0.0486781190529994, 0.0743146526156907, 0.554198559589315, 
    0.165702885592698, 0.140298799544904, -0.309144919532918, 
    0.113690304236558, 0.516976197336114, 0.48506396894497, 
    0.290894931091538, -0.100769965549795, 0.515522807611575, 
    0.268802950673175, 0.0554571841673488, -0.0355961843892338, 
    0.218827985674793, -0.0317326577865422, -0.29402524365599, 
    -0.226435109897015, 0.204620051553037, 0.367777874218707, 
    0.150341055203261, -0.176143414491996, 0.145649504703489, 
    0.0259154276303086, 0.0273262047353615, -0.460258825047427, 
    0.000949333454591805, -0.271813404488956, -0.321068490899728, 
    0.182755037597578, -0.396109056718505, -0.0686928683351635, 
    0.0413760269999881, 0.103253574165202, 0.147723925456333, 
    0.158505799203158, 0.151600414034714, 0.19432863911719, 
    0.191560709547601, 0.0860366892370671, -0.00956718785531444, 
    0.498583721186881, 0.245012585269119, -0.034501286321922, 
    0.0193800708663712, 0.634793205630839, 0.213545547746712, 
    0.109585244817699, -0.110828623100252, 0.473823745823827, 
    0.278818492262482, -0.00916634464499579, 0.00331182351399564, 
    0.608256473638789, 0.363062922183757, 0.113994213101483, 
    -0.106639645276913, 0.0868847299724058, 0.0782751424415191, 
    0.849864099803031, -0.116169741328992, -0.286412120590586, 
    -0.0640135039679957, -0.226918021803725, -0.0968817438329853, 
    -0.105134883186714, -0.178233947233873, -0.128527364074721, 
    -0.183596061490788, -0.188175545605515, -0.160520044340127, 
    0.0144642328190529, -0.111234940714919, 0.0230382231034231, 
    0.0081881694613002, 0.051810222865906, -0.0690438213959633, 
    0.00416272661712867, 0.0277267300870506, 0.127565781364616, 
    -0.0440112286020662, 0.181779897488975, 0.124903836940119, 
    0.0335181252664025, -0.00128351394739172, 0.311158260485626, 
    0.123144907716511, 0.0560450873310256, -0.00339762955101547, 
    0.164603541894123, 0.0566450844663369, 0.189014392934135, 
    0.695321618563956, 0.309484026585002, -0.236487156677186, 
    -0.0687489715515498, 0.756339669331895, 0.39889230002731, 
    0.148729570570196, 0.805127413320372, 0.319394317997846, 
    -0.0551896282049704, 0.0101495352518969, -0.168722403654917, 
    0.269811679765856, 0.165094651227808, 0.12188543414639, 
    0.115892939235267, 0.0610647111245657, 0.329994368218125, 
    -0.121483214802925, -0.203210321679937, -0.0761303021849405, 
    -0.13153467665519, 0.0114701187540153, -0.0454437279778613, 
    -0.0343619250860413, -0.0935200032458026, -0.108528694390779, 
    -0.130769309935302, 0.0726206043002459, -0.0907439143383429, 
    0.0989298413226485, -0.141174616224941, 0.022943981527302, 
    -0.162197091527366, -0.0847051912343699, 0.0199801338825812, 
    -0.0822198035307439, 0.0930349967890848, -0.0900593521967218, 
    0.0540877812035122, 0.0491009934880687, 0.0552418495724181, 
    0.0303941036916757, 0.0230729951626053, 0.038094573490743, 
    0.0566520305486397, 0.068727699354443, 0.0698896195213867, 
    0.0161448259635759, 0.028817034838902, 0.0286775464980239, 
    0.240157685966509, 0.293920215588078, 0.148013838885305, 
    0.00764199434252166, 0.308767861298416, 0.208481162212995, 
    0.161648626365085, 0.270193061929093, -0.067182562817848, 
    0.467280108148698, 0.304022531411869, 0.17878095898775, 
    0.765707793636241, 0.632080653840845, 0.141601033746244, 
    -0.230144457349554, 0.241814831280376, 0.521599416315596, 
    -0.204256240069582, 0.0505775292816357, -0.232647119359787, 
    -0.0716055855865075, -0.147213377307542, -0.0315924535320473, 
    -0.130736629762902, 0.0363279062759701, -0.205325891701753, 
    -0.0457171345899781, 0.0117322254119472, 0.0342329122890047, 
    0.0887516434742841, 0.0848441615192056, 0.143534348014479, 
    0.0828673900449794, 0.0995470853757774, 0.124697628618123, 
    0.0929207885112981, 0.0274859751199744, 0.0451964166692183, 
    0.132476196047519, 0.122361424738283, 0.0839609924601693, 
    0.0827039984942102, 0.154799475459268, 0.298613911022754, 
    0.110042731320184, -0.15490687965606, 0.0208152159029766, 
    0.497181396667053, 0.0217747982216398, -0.133490150084586, 
    0.139940016376302, -0.13727999213925, 0.920615006892906, 
    0.376591456912338, -0.126838375107641, 0.577512210106539, 
    0.437089013995982, -0.338042218183167, -0.0662264296291484, 
    -0.0884709175846879, -0.0894224767248532, 0.0147502826603846, 
    -0.112237299388851, 0.0772584232222373, -0.222104425055873, 
    0.00696019642396226, -0.0873022430588961, 0.0160901081849526, 
    -0.107796194231084, 0.101596624667507, -0.113028361956567, 
    0.0974782660162026, -0.24455025637001, 0.0473303627347465, 
    -0.140818475782555, 0.0313301819383021, -0.280442123979234, 
    -0.0495581355684496, 0.0228793988115334, 0.0604826311696136, 
    0.0714937100017167, 0.0640912724255244, 0.0791950869537147, 
    0.121277529442361, 0.143516323040083, 0.088846252367077, 
    -0.160499643734615, 0.17346447528903, 0.358044548648171, 
    0.129679821950502, -0.0286127512375564, 0.569249240774088, 
    0.288261821111871, 0.100950668002781, 0.0563144010302038, 
    0.0682754603634345, -0.00924696804543065, -0.0971777571594964, 
    0.839032976563194, 0.596207412367662, 0.171389153536254, 
    -0.619954643196492, 0.365677440601702, 0.402796199210314, 
    -0.0623569782870688, -0.0434546715085562, 0.222009672074488, 
    -0.320421055131563, -0.192680632447713, 0.0160410622815141, 
    -0.207087894473704, 0.105051904252947, -0.161412244470443, 
    0.0632619697373608, -0.0888350119393637, 0.0788478476620403, 
    -0.228614221325936, 0.0108911570647364, 0.111565877527606, 
    0.162864755126904, 0.20436738733349, 0.21140089795901, 0.166428949310057, 
    0.159655049207396, 0.232078712737946, 0.232525952566615, 
    0.160975552121927, 0.134013940938003, 0.170320906265305, 
    0.24682909882913, 0.229484276951891, 0.14551336570861, 0.148942960781266, 
    0.330199161586348, 0.242616360069214, 0.0338638955674823, 
    0.0270778553700551, 0.659877918679681, 0.25103722133529, 
    -0.132252932415497, 0.420529384446774, 0.287818330460832, 
    -0.0631301071805328, 0.0859351728659753, -0.544812154218915, 
    0.470549026184696, 0.478541470009138, 0.0926742162999205, 
    0.0222635949893076, 0.073296084887615, 0.204356687409859, 
    0.262907785259491, 0.249244170954136, 0.2016590054661, 0.149504914229025, 
    0.150774552382843, 0.211169381358719, 0.210046021412707, 0.1582616682137, 
    0.122885984996637, 0.155499796068064, 0.178437122461802, 
    0.115844602531133, 0.0617938294309285, 0.130540188545811, 
    0.183186635596864, 0.205977364983921, 0.182629659843969, 
    0.0230156585509265, -0.147963017733181, 0.177001746844918, 
    0.465518117048248, 0.258295543695421, 0.144543323794385, 
    0.157153910200115, -0.0373781093847542, 0.61313594924504, 
    0.165553221533334, -0.0033006321490899, -0.123818091698166, 
    -0.0817567578842539, 0.508184171918592, 0.0988834194291505, 
    0.0995828432332926, -0.172147379877895, 0.413880602293319, 
    0.128135734421817, -0.0882967133695234, -0.01706365779422, 
    -0.264457182570875, -0.0935783804499609, -0.279937397160156, 
    -0.246889755530385, 0.0863756280855526, -0.084122821623719, 
    0.154886488914945, -0.193230148812951,
  0.0572736678033119, -0.0536811791642671, 0.112534754796535, 
    0.00631068533297526, 0.105587851154265, -0.146378234061715, 
    0.0314142275857215, -0.024386423893037, 0.0507390640148747, 
    -0.271291298627987, -0.00876953354777021, 0.0735924028993977, 
    0.0661221393788597, 0.0831642695682056, 0.0713640694552445, 
    0.077103615715586, 0.130253856020599, 0.110140614447875, 
    0.0528756054135679, 0.0700463567320704, 0.125903599371475, 
    0.129212556959369, 0.138916939539754, 0.168984181539807, 
    0.172646810276973, 0.116277784754063, 0.0998924246725208, 
    0.199913639525728, 0.12487591982268, 0.0864409697706989, 
    0.233058916636709, 0.50035244159336, 0.411730406018286, 
    -0.226097757232467, -0.473019184850228, 0.390064287296843, 
    -0.285242141268489, 0.246255796580911, 0.495414138713276, 
    -0.0174356212411612, -0.277644481059498, -0.116154229511758, 
    -0.0264977534169845, -0.16188361823548, 0.029083787045237, 
    -0.231807032889207, -0.0247565947875573, -0.17347324853443, 
    -0.101662075215508, -0.0844045161745859, -0.026229082682627, 
    0.0491198838421366, 0.0667614014337764, 0.0791341343821629, 
    -0.00714420194722476, 0.00786764141944314, 0.100430503182877, 
    0.0988591317953953, 0.0365158867529199, 0.0901179280672782, 
    -0.0968740756701629, -0.0416290440731506, -0.00301099127196831, 
    -0.0564876234924661, -0.00571699895556144, -0.0414107546052374, 
    -0.00202474016843328, 0.00807998668637497, 0.113329008339802, 
    -0.0838898374695892, 0.0508602742493509, 0.159497577725126, 
    0.279758887740296, 0.185702776173257, -0.00131694464712749, 
    0.0976472106270846, 0.308122938528593, 0.441202645753163, 
    -0.0722300600938997, -0.159663041244956, -0.485698712441373, 
    0.236370895151737, 0.71950128104569, 0.155919277660323, 
    -0.105655457400499, 0.18675095032119, -0.173587422104993, 
    0.358000861370505, 1.1153592519865, 0.0202151438225281, 
    -0.278881441958685, 0.0122284260316171, 0.502815751798526, 
    0.0768749605446917, 0.05244989618599, -0.139469142826075, 
    -0.0681498595165698, 0.3714286429528, 0.33768892281583, 
    0.0173041525133639, -0.143814516736763, -0.108215653237179, 
    0.1646233504606, 0.114025145058435, 0.078641231314334, 
    -0.0848165981585121, 0.140240922757316, 0.0638418167023172, 
    -0.00233286225230173, -0.125906261174873, -0.00749628749532634, 
    0.202628702054844, 0.105559120050041, 0.13386387289995, 
    0.294974652836565, 0.16580103978457, 0.161026068181486, 
    0.276003397980801, 0.016607825957155, -0.111857376197492, 
    -0.159943235574134, -0.0160470176514332, -0.148716842486605, 
    -0.128341277457474, 0.106324136200135, -0.142041453074162, 
    0.0254405582355718, -0.0279760166667069, 0.0488311641207003, 
    -0.184514265058117, 0.0191892520458763, 0.11903349840521, 
    -0.00934848176671495, 0.175370044105297, 0.231988739860843, 
    0.0838860102189576, -0.0371949648980737, 0.113818204337819, 
    0.311448819755471, 0.251489692422608, -0.233682571458838, 
    0.53856296738358, 0.502702205139206, 0.205018814973675, 
    -0.280621788388243, 0.904462896813003, 0.451033704710135, 
    0.204770617143467, -0.28571758689643, 0.524108363929431, 
    0.377818971993125, -0.0284021426464259, -0.00689160465758516, 
    -0.215694054515982, 0.163065810499249, 0.252511514823627, 
    0.0822066023756493, 0.0227913655880542, 0.0143583045098165, 
    0.259027521529834, -0.20429916257696, -0.196501292552544, 
    -0.166504440769859, -0.202614131670448, -0.112338202032802, 
    -0.21998388818732, -0.132959302851514, -0.160301838289964, 
    -0.000641424968124971, -0.217933820396817, 0.0478281565615012, 
    0.0577272481330525, 0.0969644144316465, 0.013364750354693, 
    0.079468360869285, -0.00441020273498109, 0.0512289753396796, 
    0.00397072240079967, 0.0469242810223485, 0.0451835333068275, 
    0.0664308518598461, -0.0115456966312015, 0.0322658245051752, 
    0.0191464358989268, 0.0420729570135327, 0.00487167186822618, 
    0.040942740212313, 0.0125952941166855, 0.0384041445837405, 
    -0.0275998671792894, 0.058146580031036, 0.0490390060217512, 
    0.0841434569382775, 0.23161864833997, 0.139135113898871, 
    -0.00475080794584448, 0.042869723494974, 0.357408016415769, 
    0.129920316428167, -0.278572967856206, 0.25497954501914, 
    0.409301404022097, 0.109900679982411, -0.381134160417564, 
    0.117014235094782, 0.794692728419421, 0.319049257325814, 
    -0.0697771647841968, 0.212270408337388, 0.538736663213336, 
    0.184336329475732, 0.118114306641846, 0.0369396175759994, 
    -0.164612106661607, -0.037292774754356, 0.633221829442956, 
    0.0694298530646156, -0.210666539134465, -0.24070567996129, 
    -0.136507092530822, -0.0723506050711822, -0.262723037107912, 
    0.227155218463003, -0.240289125086871, 0.14608835392565, 
    -0.180249466462659, 0.0413525167594666, -0.101433743196036, 
    0.0822727718369237, -0.320474903127973, 0.0261941497297721, 
    0.0469240965464819, 0.0614124099087221, 0.0867602592729415, 
    0.0842757180759558, 0.0711465200865887, 0.0878951799241905, 
    0.0484889669945775, 0.0812959664340954, -0.0141577447178988, 
    0.0739022574399402, 0.137666685872984, 0.343065341941476, 
    0.233940346291985, 0.027459451186088, 0.0621532556351512, 
    0.427699748561315, 0.266172886554916, -0.0238938769731793, 
    0.272877888043781, 0.597351496566931, 0.0990597353495892, 
    0.599525614356828, 0.57963263475499, 0.0641593074141628, 
    -0.00300095571996251, -0.137731188605062, 0.547560098406961, 
    0.757832683805442, -0.305131957364501, -0.246450794429203, 
    -0.0909583041221123, -0.141962719388661, -0.090590311412845, 
    -0.155033428915618, -0.0497741854310935, -0.197014583988981, 
    -0.0618097499630367, -0.136643384363348, -0.141145740832259, 
    0.0247944987510734, 0.101283687809689, 0.0904387929876464, 
    0.113857962918936, 0.0868805265621897, 0.103613272331525, 
    0.083517581941604, 0.0875982441526417, 0.101386619526459, 
    0.0884805280075826, 0.0951438159098306, 0.10605435059623, 
    0.107254784456518, 0.114953289751204, 0.132234499427472, 
    0.114118168968263, 0.115888679178473, 0.162351436990382, 
    0.123346494502808, 0.0107886508064875, 0.235488259388764, 
    0.227434157897807, 0.0502213482976991, 0.294257078394645, 
    0.314718537249498, 0.0915302033229291, 0.308428914323026, 
    0.397703550757061, 0.0805578379006992, -0.00719218985612199, 
    0.387990079935416, 0.429921838351688, 0.484534257731704, 
    0.310004996680315, -0.203764061946725, 0.792508075070954, 
    0.443836848531719, 0.0639868929262964, 0.658977251874264, 
    0.326763672310485, -0.25011588593051, -0.039517205995205, 
    -0.160677105136087, -0.0655409769225084, -0.136827916192134, 
    -0.124813518842682, -0.0971120574125759, -0.0202007080742902, 
    -0.151216379888304, -0.0360377734035495, -0.0332387653741425, 
    0.0219569654306971, -0.158999195675803, -0.0514890780431885, 
    -0.0172342370989507, -0.0104773095333365, -0.180202375589227, 
    -0.0390309042843945, -0.102178587522574, -0.212063429871548, 
    0.0324544826427688, 0.0520997799116661, -0.000569819194505231, 
    0.105826331756198, 0.078526529909868, 0.0823927300322767, 
    0.228555700918505, 0.0751529560363278, -0.0319011649418702, 
    0.228320537517769, 0.190157268605765, -0.329287525597475, 
    0.00282409111166358, 0.731123627012608, 0.385075312480938, 
    0.168774804931689, -0.341434236243023, 0.0332280149702709, 
    0.530806324341885, 0.282238220571788, 0.0546828070647791, 
    0.149776058645505, 0.11597663111026, 0.0365013107321284, 
    -0.0244265753245877, 0.109391127510717, -0.0217770277747059, 
    -0.0556586677541351, 0.0396822199012802, -0.0272639975529114,
  0.265600326779809, 0.317981917863409, -0.344681343507994, 
    0.421173424442961, 0.670691745479535, -0.452269816209094, 
    -0.39737142850589, 0.103118278997469, 0.852151101027247, 
    -0.327388840171752, -0.0869659041797881, -0.116325526893117, 
    -0.0435850933431622, -0.161081285537695, -0.0607228134147605, 
    -0.127978290247012, -0.106712253485454, -0.110709805840253, 
    -0.0962095738417141, -0.117867009654275, 0.0157801702039565, 
    0.00919659743677076, 0.0509086211808406, 0.109288369514609, 
    0.0868744549349527, -0.0476187763660653, 0.0914410851740816, 
    -0.00718311444886807, 0.0526921796603447, -0.0296793860448199, 
    0.0257727843808408, 0.0714889190238626, 0.0894586415767948, 
    0.0812590999239891, 0.0823065120356192, 0.0777750504942932, 
    0.0922812644675727, 0.0997055345577802, 0.0241226346591014, 
    0.11983251390417, 0.300880595354316, 0.10355863211042, 
    -0.00885196523003291, 0.468548014428129, 0.246941341080973, 
    0.0939021495762441, -0.0386304521534842, 0.22910902109563, 
    0.291484681153869, 0.394924776619516, 0.277321256091122, 
    -0.0440878314341743, 0.452156111578883, 0.552998246241855, 
    0.228634576871646, 0.251798156449412, 0.610100525072789, 
    0.0183223219316704, -0.0557404654695584, 0.0919792591534953, 
    -0.268112270368787, -0.242677641760712, 0.158505411820023, 
    -0.265050162348293, 0.0370772311883169, -0.0516690733662894, 
    0.0826920960918385, -0.160623305972524, 0.0971726979190612, 
    -0.153863859498259, 0.187678977611932, 0.1197266716922, 
    0.147968715181559, 0.129879152010781, 0.0590831958172783, 
    0.098291502219162, 0.172664071358501, 0.156266104039541, 
    0.0950759843423239, 0.124735627206895, 0.105553944133401, 
    0.105005420312204, 0.126657730155273, 0.126144330467471, 
    0.112586065780864, 0.11629270915726, 0.110929479135056, 
    0.129175864141559, 0.131175445928212, 0.109200919224795, 
    0.106005374936807, 0.0299081191268474, 0.231412677720331, 
    0.302269973158891, 0.166956047556899, 0.0779254061108372, 
    -0.030995416387833, 0.30868514519773, 0.371986032934905, 
    0.138137422422506, 0.0484549528743749, 0.254831923915569, 
    0.539744514923281, 0.0232675493421884, 0.52873179076706, 
    0.507325979406506, 0.435523102970757, 0.936163348679887, 
    0.303122063478536, -0.134526461447724, -0.160978138750903, 
    -0.182425183710111, -0.133933202574153, -0.145308726998088, 
    -0.196690337322813, -0.0695552220900431, -0.202751884384497, 
    -0.0808915887809401, -0.176044295250335, -0.105232339049681, 
    -0.00687172886937169, 0.0191653491186067, -0.0199898107230772, 
    0.0076923736351537, 0.0403177320224395, 0.0593671930968418, 
    -0.0295244687026882, 0.0547982342141144, -0.132132756993655, 
    -0.058262307412233, 0.0104934033831754, 0.022547782782811, 
    0.0335506903904975, 0.0388782468756118, 0.0366853545441357, 
    0.0322010677342418, 0.0191644360130976, 0.139678285431902, 
    0.235809183684266, -0.238516742560135, 0.394374292884466, 
    0.289516831382768, -0.126748209686824, 0.242657363692294, 
    0.591416916494975, 0.147725507105926, -0.088906556025042, 
    -0.0650502013142013, 0.691557565754081, 0.356887499839751, 
    -0.120602791544883, 0.777149929591419, 0.333343599840366, 
    -0.185834702073126, 0.310889012167844, 0.562240130005485, 
    -0.0036019109395261, 0.499408405635994, 0.632356378753863, 
    0.0342705742508426, -0.0460870214518522, -0.0076787233332475, 
    -0.026720987818906, -0.00321301710360733, -0.0179942380432326, 
    0.0596500542433108, -0.0582662107404086, 0.0413031298773114, 
    -0.00319678473436652, -0.0662740390888169, 0.351329055653669, 
    -0.174895069116708, 0.353060054702878, 0.609389242511327, 
    0.145649891033588, 0.0270857250687508, -0.222541049787811, 
    0.0258192929901822, 0.609712758513708, 0.219261388662446, 
    -0.0174742168014712, 0.105595428900514, 0.72952830308932, 
    -0.0654288978944116, -0.368612130092388, -0.0711080895947178, 
    0.776749801783802, -0.0224403321628886, -0.125305014987418, 
    -0.119514569716246, 0.618585645719245, 0.219241961630218, 
    0.0311832807000558, 0.138330513470755, 0.227047523397654, 
    0.110794505501682, 0.445852766999239, 0.449838843410916, 
    0.338620663425732, 0.678144106387067, 0.248918679837862, 
    -0.441326473347878, 0.0593820944737826, 0.735823766471807, 
    -0.00135620052512028, -0.174380045286546, 0.198782778784356, 
    0.0198652736090935, 0.176325955812618, 0.884343659110352, 
    0.331917027640925, 0.121938936756602, 0.13633455549998, 
    -0.191078474709706, 0.239007386543335, 0.165203720253471, 
    0.00035830767845435, 0.569331585852792, 0.278257315627143, 
    0.000921542267104364, -0.110060809345407, 0.0871945146565885, 
    -0.090913394968047, -0.0550074451107095, -0.15134373382839, 
    -0.133367142790457, -0.0637166099184538, -0.148500474165152, 
    -0.070549869925819, -0.100560171613241, 0.0771788228476892, 
    0.0818655652010852, 0.150493034865522, 0.127038758943274, 
    0.0838594880252107, 0.0639553845897003, 0.0793847164789562, 
    0.168844939590165, 0.126633149512942, 0.0568566857214311, 
    -0.0311237125487798, -0.0123467553463744, 0.0556682159330953, 
    0.0173802168673182, 0.0749598663725484, 0.025694776772972, 
    0.0576300361986018, 0.0420917771450459, 0.0581698738113496, 
    -0.0246274724264188, 0.0417291003554351, 0.104553575043294, 
    0.0840151391670415, 0.0672654728900737, 0.181930816391627, 
    0.198866486160401, 0.113355712218037, -0.0750404567545145, 
    0.303862993877658, 0.23030137170643, 0.124525843982284, 
    -0.148356656057903, -0.0649807267460477, 0.498525765392471, 
    0.474065067453113, 0.469053802019042, 0.418160032399553, 
    -0.0990737030272392, 0.740027194517871, 0.734545972982207, 
    0.349376212634525, 0.156488560694749, -0.186364761311433, 
    -0.0744835091350079, 0.340840343285273, 0.104454033909186, 
    -0.0779598912409238, 0.240682580464105, 0.0950591706784597, 
    -0.141086601509361, -0.170003639128992, 0.120338278379645, 
    -0.253347688733543, 0.0356744451156539, -0.324521167111101, 
    -0.14185608471637, -0.0974638436502712, -0.180375550905095, 
    0.00342901270160025, -0.152759395305328, 0.255118255691126, 
    -0.00182596258005681, -0.0260579336482496, 0.287325634106171, 
    0.416666257954321, 0.148352989800247, -0.358818937726536, 
    0.304942007172906, 0.474970014823517, -0.373027433369495, 
    0.177229175229499, 0.85065749386875, 0.13295527853862, 
    0.0758050265658018, -0.312431038021377, -0.0214163529718602, 
    0.469841012296489, 0.740809404059665, 0.611716278176595, 
    0.210379604445121, -0.232865477066461, 0.299177079463585, 
    0.324526976407936, 0.0835008186751163, -0.00684109384192785, 
    -0.0930211791699718, -0.0474456739546963, 0.134143828617646, 
    0.0248582537649285, -0.0429630376828921, 0.159304114737652, 
    0.143120629944623, 0.0918366127684027, 0.0639126796755139, 
    0.0757698089380857, 0.149482136326475, 0.0139230930186121, 
    -0.00898415658466362, 0.023719931542682, 0.104702488340164, 
    0.0466464527864652, 0.0361464605119274, 0.0473516460312653, 
    0.0545329613762218, 0.0581308331203844, 0.0498789642444357, 
    0.0451701257429067, 0.0683728341649606, 0.045769153445932, 
    0.0431203335032567, 0.0433966732072225, 0.015593510994761, 
    0.0502368445445521, 0.0296560398092379, 0.0438343090191224, 
    0.0376310785471191, 0.0597781157006808, 0.0332609445954721, 
    0.0712555868752043, 0.00488954978611918, 0.165046425185224, 
    0.112904076511902, 0.0544492415149118, 0.320299754814275, 
    0.171428422887601, 0.00531865659887334, 0.144758866347828, 
    0.289099261087161, 0.0319115696477868, -0.127332293157817,
  0.176588157100965, 0.152154823265459, 0.143678097070958, 0.239346425087059, 
    0.282413380721278, 0.217173132126632, 0.198137989007952, 
    0.265106372133373, 0.23103527575426, 0.191749583603471, 
    0.348611565881787, 0.339489240890788, 0.141897088021361, 
    -0.00335457676006508, 0.484681130893413, 0.319229965602557, 
    0.0710109779869723, -0.145628640002381, 0.379537053305866, 
    0.454517136905473, 0.182771052713238, 0.0106639913776851, 
    0.165011345160865, -0.0588978600399128, 0.190152324657859, 
    0.753797167529565, 0.408749893609891, 0.0751947051206068, 
    -0.410565922120447, 0.019867811285691, 0.568403017338331, 
    0.136714926225204, -0.0634862635606418, 0.271988546541591, 
    0.249892004749858, 0.00105187195248187, -0.379039209985118, 
    -0.00040634583980137, 0.312959836431388, 0.144248657231118, 
    -0.0757121015355392, 0.0904287765002012, -0.175903324892621, 
    0.0274342037795381, -0.221450306489978, -0.0540573416354156, 
    -0.164295816546091, -0.137128790621441, -0.0286553403958193, 
    -0.161816002039922, 0.00806938278382739, 0.0920492391539024, 
    0.11356085839185, 0.168101672491848, 0.229593937070196, 
    0.157459103988573, 0.097263142863844, 0.280205944412454, 
    0.317143831241048, 0.225429825321163, 0.189125222505222, 
    0.0303920603607941, -0.0741652940900105, -0.0341820256637552, 
    0.84256852589665, 0.33372782191122, -0.0870003749821897, 
    0.387910109246109, 0.498221606482519, 0.0997372954273977, 
    -0.0826787110236915, -0.0233731650718292, 0.83033803802159, 
    0.30644968199693, -0.000828598140344153, -0.195748582007901, 
    0.206475993567466, 0.664685546801119, 0.333786293023396, 
    0.0890170573357197, -0.131045991231581, 0.246953570194001, 
    0.312660293744186, 0.192576062233394, -0.0425779078040717, 
    0.322257186921021, 0.0567857248861829, -0.0831603574475971, 
    0.233841517319357, 0.0191088780561767, -0.152985437860799, 
    -0.0527524131392059, -0.168175106617058, -0.0779629246593729, 
    -0.0536987507553434, -0.0996307563990213, -0.00394664285440024, 
    -0.191395957073356, -0.0206687389782856, -0.114815662596583, 
    0.07510049421377, -0.109907015282683, 0.0216369370566201, 
    -0.034128270970872, 0.0370308191785056, -0.0730448598686431, 
    0.0439299554879038, -0.0531836817113113, 0.0448975369729852, 
    -0.129194030122423, 0.0566452502452142, 0.0197111911582831, 
    0.0634459894632814, 0.244648918254815, 0.137960671211443, 
    -0.0313925387154652, 0.0566557640992048, 0.464874164760863, 
    0.194972183697097, -0.385700218359628, 0.258587765527051, 
    0.58896948327293, -0.027952452887986, -0.0512898896438779, 
    -0.207050332030145, 0.598466563707874, 0.137876582681504, 
    -0.138582647832062, 0.370259203739568, 0.491431192503052, 
    -0.194470004535928, -0.0502317531517766, -0.0441266059097528, 
    -0.0626776654812389, -0.0612470157130711, 0.140085797617178, 
    -0.194367404709901, -0.11668410152357, -0.00244175634903249, 
    -0.0165153402355293, 0.13154079368077, -0.150351440165651, 
    0.0952732973093299, -0.0070976631494728, 0.0780676198387533, 
    -0.230064805363023, 0.0383993682116213, -0.126403711437949, 
    0.0290608861257187, -0.313545077184048, -0.027398293068944, 
    0.0453057766030357, 0.049630750120507, 0.100217756587436, 
    0.13577697915446, 0.112773977577995, 0.133433467484414, 
    0.184396276507027, 0.119114933110975, 0.0383319945387022, 
    0.0987204421013625, 0.023632661434143, 0.214100731247632, 
    0.525425409271958, 0.267939471399964, 0.0849711174819761, 
    0.599331503368353, 0.206615692123251, -0.053029293905799, 
    -0.121683623612514, 0.784697296766675, 0.108548202918234, 
    -0.185351472658623, 0.0599773049785086, 0.631527521526282, 
    0.608725989902903, 0.335482931881329, 0.0745620509756178, 
    -0.41475858012273, 0.0548596677704212, 0.402820003840785, 
    -0.141681803779414, -0.198295440712073, -0.0500542129435026, 
    -0.236556000237268, 0.0695910889978251, -0.244748592648973, 
    0.0168001772681895, -0.248593720071971, 0.00618476025554878, 
    -0.0290497859675744, 0.0945184684263655, 0.0403180932695746, 
    0.10137599804099, 0.0295466332699216, 0.0850017043799105, 
    -0.13328295463152, 0.0251343060044723, -0.12130530884184, 
    -0.0849291284605208, -0.00281478096705927, 0.0638133395325847, 
    0.0278340685150877, 0.0490349550658862, 0.0438653090400394, 
    0.025002752457483, 0.034461321833102, 0.0689396265387663, 
    0.0630619815495547, -0.000691672093171031, 0.105523501643821, 
    0.137493896581043, 0.100094166537759, 0.213859682677491, 
    0.266648524781617, 0.122555575777718, 0.0835526430761312, 
    0.379925621536444, 0.213833962217663, -0.0439639164253157, 
    0.410952902090198, 0.385507237112117, 0.0564162713351136, 
    0.652213736504179, 0.435639839521556, 0.0931298431522912, 
    0.0870010602098521, -0.327292507939657, -0.152525440004884, 
    0.500050687553638, 0.44517710056282, 0.186237699171104, 
    -0.0321039725872626, 0.310081749293849, 0.217478976401722, 
    -0.13700507398264, -0.435311385336852, -0.13410943388385, 
    0.496491630028764, -0.000820377587322521, -0.140184841647982, 
    -0.19817283448606, 0.0287172072417371, -0.0897464572524607, 
    0.0487078111536948, -0.278248898840177, 0.0275087882557914, 
    -0.153229273648165, 0.0132269276320938, -0.299695081405713, 
    -0.0547070826264651, 0.111201877693745, 0.10636055684947, 
    0.10498771278678, 0.220847561029646, 0.248004919666637, 
    0.222991394031199, 0.240203120330583, 0.187179841822182, 
    0.128467987268562, 0.358439372189798, 0.351400819119822, 
    0.141270359816536, 0.248825659129606, 0.610070136365626, 
    0.287528888704366, -0.0722596950548925, 0.335986054964361, 
    0.646197269143534, 0.214219100831364, -0.0907529306145367, 
    0.507711289652607, 0.35497748330582, 0.0415208382453126, 
    0.511283901293774, 0.447516042441014, 0.078644255392938, 
    -0.228151728465384, 0.425756171261755, 0.56332302700549, 
    0.0106867151184415, -0.113137421684581, -0.113064760170483, 
    0.413286663214324, 0.144581690264819, 0.0488919163888816, 
    0.0618418330671629, 0.00224348020545953, 0.00974438309478043, 
    0.552002870287224, 0.173809354548586, -0.00437057251219455, 
    -0.0108404732978451, -0.0190790865744266, 0.0163126833529032, 
    0.0229255081217602, 0.187396393278701, -0.0474572083108528, 
    -0.0507913381128763, -0.0564644211780889, -0.027957717224651, 
    -0.0816925540673161, 0.0920422614916151, -0.153386185142602, 
    0.0186340244981841, -0.0965959509958757, -0.00341621061591613, 
    -0.0483825566787852, 0.0427797107047647, -0.156886345803295, 
    0.025184557552736, 0.0711931141098906, 0.102808657328602, 
    0.149427003622301, 0.117547023953681, 0.152075968220665, 
    0.449895424453077, 0.235112125615582, -0.18926717132727, 
    0.282392730216604, 0.484007495066179, 0.141651516038866, 
    -0.335263484229943, 0.30196531083448, 0.641284692960443, 
    0.0676436351316261, -0.0751858158360129, -0.111217384414881, 
    0.641137044825758, 0.0172215394102153, -0.13008813885567, 
    -0.0826015107944886, 0.0664326831319939, 0.117826849205302, 
    0.288818704714014, -0.0160178199593299, -0.133581036050204, 
    -0.119277170015803, 0.0315831010904928, -0.0511317195670615, 
    -0.0719160070640131, -0.243051474183166, 0.213637421118577, 
    -0.28386111961551, 0.0849420412507149, -0.361802894782862, 
    -0.0419727829304162, -0.122850331974335, 0.084581813078971, 
    -0.488294124107904, -0.0154077123358132, 0.074640578326536, 
    0.014685579932305, 0.16995584549449, 0.216469617520026, 
    0.124296860536803, 0.0983258589638733, 0.174122579289935, 
    0.168289764258217, 0.123640607510391,
  0.0947021049875212, 0.0261552932998275, 0.107774779263539, 
    0.0129503739576857, 0.0629584365874055, 0.026767195815874, 
    0.0450284819277309, 0.0576363539668189, 0.00365589667865607, 
    0.108312218990733, 0.4476341350577, -0.277874045810742, 
    0.306805836817598, 0.620347921993004, 0.153014811610928, 
    -0.0331074473802989, -0.124930721624561, -0.209872700173584, 
    0.536731347549741, 0.47874916161694, 0.169573722505407, 
    0.150151816418625, 0.293077178563487, 0.102009682476491, 
    -0.121234120335493, 0.780353090946909, 0.265976120944928, 
    0.0733900169021862, -0.128819390851476, 0.566484567317412, 
    0.211256689247219, 0.0526461786830727, 0.03140610439607, 
    0.0593745919255281, 0.0667862849225085, 0.0430923507836755, 
    0.0311091551339184, 0.0813965583576907, 0.11077761351534, 
    -0.166857162552486, 0.322725696210897, 0.287964048580162, 
    0.140900270271871, -0.203585088555507, 0.640953594823663, 
    0.223004698901115, -0.137915427706005, 0.412607421181446, 
    0.295009761444906, -0.0225394434544144, -0.194963408196678, 
    0.395957899385011, 0.554491774644292, 0.0906743273331455, 
    0.0723587707425443, -0.57523219326696, 0.459725304295563, 
    0.425629927075933, -0.227375584871375, -0.0240198612402099, 
    -0.418816166293717, 0.0399158928510687, -0.312998696160181, 
    -0.211762739326804, -0.0339083699981337, -0.205872658751817, 
    0.110329224217063, -0.160532136730733, 0.118291930329959, 
    -0.138390473105091, 0.143016938663397, 0.0259855688415507, 
    0.0662988416086, 0.0343403121148106, 0.0725198951945147, 
    0.0581579220728179, 0.0925828927546997, 0.090903277613749, 
    0.058649799224365, -0.0575490080148847, 0.0180762588563027, 
    0.0457462973966983, 0.0520197132784584, 0.0644049751981477, 
    0.0708215599965001, 0.0553807727986797, 0.0637244103741643, 
    0.110787986034333, 0.0246879078139655, -0.0555728460780196, 
    -0.263456002497459, 0.417776496139672, 0.339307432311888, 
    -0.0145894310652784, 0.35204768061642, 0.502038101242766, 
    0.191594344809344, 0.0627690550823956, -0.069515298082018, 
    0.619500615597947, 0.236079855541927, -0.0161908096903528, 
    0.247502561255339, -0.545169064669842, 0.233192112011423, 
    0.369118897199898, 0.497472431613128, 0.365739051041135, 
    -0.073358770783605, -0.0398547330260658, -0.375189702385757, 
    -0.0903068107535667, -0.310724927971063, -0.082144693382227, 
    -0.303330266673343, -0.174670955970206, -0.0554785073463793, 
    -0.215958045936517, 0.0983041783668616, -0.30121568351478, 
    -0.0180100808396612, 0.0568093194960722, 0.125166282848875, 
    0.195692269627049, 0.240069632752275, 0.223576217420004, 
    0.203154833072053, 0.216392908769468, 0.220143616715027, 
    0.205618978400572, 0.233808244511419, 0.214563093230088, 
    0.233053675155182, 0.334166858210945, 0.319550603944373, 
    0.199514234788913, 0.170021673993399, 0.317173440889359, 
    0.362202402220627, 0.344900092246753, 0.334284577706114, 
    0.235551887008778, 0.0635580452290806, -0.182645638653179, 
    -0.209021923892516, 0.656352091884287, 0.297851064424219, 
    -0.0291699505603952, 0.327238886520889, 0.464164660299433, 
    0.434822128544317, 0.323375624097308, 0.0128233413874847, 
    -0.114001349273471, 0.0542332654992006, 0.403580313164422, 
    -0.126602995242893, 0.251970571815479, 0.438643973806839, 
    -0.011265437944039, -0.117636369758067, 0.0850244253458935, 
    -0.0932327041812992, 0.0187529748173417, -0.0322899337238302, 
    0.0601138691524996, -0.259245755095696, 0.0399428733063029, 
    -0.263571167290357, -0.160240820080223, -0.00502536056779447, 
    0.0605093965352917, 0.269896924947138, 0.207553088935608, 
    0.0524706865687853, 0.190203748017428, 0.436325329718767, 
    0.289337822957369, 0.119875606345602, 0.109602048721704, 
    0.357580412525217, 0.440437786198389, 0.350519709028975, 
    0.334690176610416, 0.388675466351118, 0.315095208926459, 
    0.181124528229956, 0.18505178022054, 0.411624866194427, 
    0.386512993815304, 0.173007507903899, 0.0282505457107018, 
    0.285503459802698, 0.431313991851771, 0.184045751131386, 
    0.0131268362816463, 0.460613577403277, 0.230491922026646, 
    -0.0151809353135781, -0.164715734790973, 0.376647712295162, 
    0.541366662749881, 0.0775525748964476, -0.228121368482318, 
    0.00789323624805069, 0.152926807943728, 0.730076981340473, 
    -0.273060941814435, -0.40402938194864, -0.0815767620017458, 
    -0.257767680934135, -0.227606244861394, -0.00602721194467599, 
    -0.259820625551463, 0.16316962147665, -0.148778712490298, 
    0.150625523021555, -0.353680859919908, 0.0265010812933086, 
    -0.153377992342848, 0.1462797389298, -0.106232223531365, 
    -0.0407708256439583, 0.0820577296350648, 0.0779705949551337, 
    -0.118878702377971, 0.0568867247113612, 0.032189465833677, 
    0.0326344246564636, -0.136617812753587, -0.00408082604647898, 
    0.0206447985336188, 0.0293608462137745, 0.0340868186756077, 
    0.0353983128613321, 0.035912089035213, 0.0317690862726496, 
    0.0237742257885581, 0.0366109158722077, -0.0105919682219718, 
    0.136385620060795, 0.0914851986068589, 0.0928696199126713, 
    0.251910552546758, 0.228832928153813, 0.154073266116663, 
    0.117093956845101, 0.205351272249679, 0.533185250382746, 
    0.100083050892144, -0.111910629884289, -0.252821438658789, 
    0.746658142641245, 0.290186576647744, 0.309657259100409, 
    0.595505451888013, -0.19882274724397, 0.78870970326515, 
    0.619374751666108, -0.143712086543582, -0.215949300779726, 
    0.122859380254962, -0.153327618505987, -0.0347978015493804, 
    0.0310298965821674, -0.0211610641403233, 0.181817794386683, 
    0.00768526347366313, -0.0804837442880463, 0.0661439579960583, 
    0.027151119224235, 0.132135588870254, -0.0310987114199326, 
    0.0925530354808162, -0.359816717959663, -0.0255554894250099, 
    -0.155435410757416, -0.206251875540873, 0.058755827641117, 
    -0.21580674397471, -0.0437573872219759, 0.143054899129282, 
    0.0876804878949974, 0.00827235329009676, 0.347070448798297, 
    0.309257228010945, 0.0986622165094542, -0.0255718875145732, 
    0.178864775622928, 0.351344338250657, 0.325080046091202, 
    0.253763353038497, 0.188588478538086, 0.175193916247395, 
    0.201768549522047, 0.203840956015256, 0.194843293154008, 
    0.199136050926242, 0.118056450314752, 0.122170874117245, 
    0.317304013872423, 0.211536881513562, 0.0734821694004216, 
    -0.0820942034196898, 0.301366382356093, 0.36382426152435, 
    0.156001906129984, 0.138381406790153, 0.451648641351579, 
    0.236463044067224, -0.102561078841428, 0.34493595645521, 
    0.320956240538064, 0.583363860419572, 0.670361378479839, 
    0.256153127678286, 0.298491434961974, 0.39299236834456, 
    -0.0635904833069108, 0.177590550232203, 0.477981263469801, 
    0.129871690769445, 0.0261674095590466, -0.173466816588578, 
    0.235149785437443, 0.257531895352901, 0.117008090453897, 
    0.04813928704079, -0.0702924663193112, 0.0285646464779158, 
    0.214205958753361, 0.151009358205849, 0.0177170589435805, 
    -0.00683656809472157, 0.146781878877693, -0.0806027530519424, 
    -0.0774016040037232, -0.0165932823438099, -0.0684139531570969, 
    0.108401821137978, -0.115261426965577, -0.0451837889999011, 
    -0.0824352286088379, -0.00831610828472147, -0.258890610587687, 
    -0.0395159413225046, -0.151228071346751, -0.193739798527486, 
    0.118900791230774, -0.246482434919952, -0.0445612868408832, 
    0.0376528853833536, 0.131769815972392, 0.148572471251375, 
    0.137660156365733, 0.104872979315806, 0.123990241553353, 
    0.181075141272326, 0.17365167338908, 0.146314810030797,
  0.14426469208008, 0.0504384433885185, 0.201841335892556, 0.366889363757095, 
    0.176221052152829, -0.0234849586855073, 0.208140615002332, 
    0.422364493034459, 0.169752167372772, -0.021023321166798, 
    0.107401958496055, 0.291880654296643, 0.688705302853655, 
    0.31500907856338, -0.287676282263874, 0.0497944720224221, 
    -0.35690734223392, -0.0041647393780061, 0.348065593749099, 
    -0.1603719585487, -0.190602414076728, -0.0671000269952509, 
    -0.160045800283245, 0.0156207444693638, -0.266507344096714, 
    -0.0372212332308675, -0.267289864540288, -0.188727112231172, 
    -0.0351626145761495, -0.14811103647419, 0.107233921425286, 
    -0.150079621587804, 0.0359049635079775, -0.0517805545388888, 
    0.0247638377599043, -0.130797343754422, -0.000468113270456649, 
    -0.0107542465429445, 0.0495265714711693, -0.138236826606916, 
    0.0127726384984249, 0.0351019618944718, 0.0383686853102424, 
    0.0357716508901676, 0.0408436308386875, 0.0265148456053595, 
    0.028420101922863, 0.0507534108461395, 0.0421542271733268, 
    0.01229636050269, 0.11580089524784, 0.0302604934280508, 
    0.0967030280981533, 0.290568522393969, 0.272286502588554, 
    0.161776564545067, 0.0715977402862178, -0.0272314406688965, 
    0.575966010170957, 0.145227094790405, -0.231729204873673, 
    0.283854391451597, 0.488920836185419, 0.0667708107656056, 
    -0.196590933848736, 0.499781324343076, 0.395207648600258, 
    0.101375712825827, 0.453310688018417, 0.582797338569438, 
    -0.0354044869297055, -0.0316338763640874, -0.0441622365346818, 
    0.0570771982813352, -0.134072679403651, 0.0505577938164326, 
    0.0627283000883665, -0.0184008544306159, 0.00682776223321141, 
    0.126324015424658, -0.0229336247967484, 0.0303710167521429, 
    -0.16555057749826, 0.00636540044342443, -0.0714183463761925, 
    0.037277833968517, -0.264994468390034, 0.0309904298904932, 
    -0.320937652683926, -0.177506599961138, -0.0300439494282804, 
    0.0346905662280692, 0.0492159907513457, 0.0783503539738246, 
    0.113838989031477, 0.0906071792308261, 0.0563989683798174, 
    0.0577697197191353, 0.0670699095787462, 0.202252309742169, 
    0.25262082145433, 0.0495253888414416, -0.229905152479583, 
    0.446525227853033, 0.36012751193708, 0.0734115580979367, 
    0.516069858885897, 0.541279757456907, 0.257781830644846, 0.2288251630962, 
    0.279011184149708, -0.351511830674361, 0.531351545714984, 
    0.456205472275122, 0.144307090444403, 0.263177498512389, 
    0.725062161629671, -0.0214137709739536, -0.474089995454762, 
    -0.144087012272481, -0.192966904094221, -0.288227395015013, 
    -0.243618863955224, -0.213859373818623, -0.258377504267672, 
    -0.209394404756056, -0.104929052943052, -0.251183773347057, 
    0.0790969994782253, -0.297495605466153, -0.0157681864540573, 
    0.114696627306487, 0.134972289254176, 0.145290074470403, 
    0.14721314221581, 0.122501447801276, 0.125379213871914, 
    0.161437096917079, 0.1617637589056, 0.0992564591101992, 
    0.103038779755141, 0.185836987071759, 0.257956404134532, 
    0.174852726081335, 0.0551940607978169, 0.14452643798287, 
    0.368022433382288, 0.307678673808023, 0.183962461456931, 
    0.143218783104267, 0.185575958988378, 0.251896242153465, 
    0.270399411652328, 0.268326868444187, 0.226762349718525, 
    0.156163245513487, 0.155010128979397, 0.252403197436119, 
    0.25238445225388, 0.231795348740098, 0.210288406847789, 
    0.0646113312911291, 0.0511446248165457, 0.525563970010359, 
    0.26867434781464, 0.0542086970960787, 0.103901044073845, 
    0.221289468226464, 0.0403049062059724, 0.592203922039946, 
    0.460070581424589, 0.111687968278564, 0.136129363541243, 
    0.243290181314317, 0.0760069621694777, 0.555522452089866, 
    0.385829173145949, 0.235733514224448, 0.876751328438733, 
    0.273166771739826, -0.143550273527632, -0.0723814429960719, 
    -0.0396788967152916, -0.153841425415563, 0.0241705712047226, 
    0.000851810488092977, -0.0260165798119884, 0.0572258881335153, 
    -0.0693454983836743, -0.104118147318114, 0.0553575335070785, 
    -0.16112717575805, 0.09734763091273, -0.0950925462821875, 
    0.0793048570403757, -0.172702223526363, 0.0620919544500236, 
    -0.113035831992378, 0.0416728378989266, -0.229378977910139, 
    -0.0348934084449439, 0.062115808012897, 0.057791481346099, 
    0.0704408054630648, 0.137126186018727, 0.146982037413947, 
    0.154827083903432, 0.154906106651738, 0.0728339603091948, 
    -0.0357511462163597, 0.488441236728889, 0.23752727177031, 
    0.0349938111953414, -0.172664174643536, 0.477631512491391, 
    0.393497304481328, 0.155368232679555, 0.0975643351199595, 
    -0.122188265186522, 0.730578804635999, 0.227641847605869, 
    0.0187795792923754, 0.0203069834037598, 0.189758902386772, 
    0.372847943323359, 0.353509151454561, -0.0514494720479899, 
    0.697010158603784, 0.446528604815823, -0.290460394936041, 
    -0.240787189968901, -0.160318673447552, -0.114857711109285, 
    -0.225007684762423, -0.095422984758938, -0.13692584173977, 
    -0.121867740581475, -0.102213522730811, -0.151490675328056, 
    -0.086366679073728, -0.118110995997012, -0.0306090954804117, 
    -0.0608503325690696, 0.0100656280575952, -0.0141864856389382, 
    0.0882383003752657, -0.353889975664241, 0.00731467452838275, 
    -0.118349742711313, -0.155950798361914, 0.0353041728016375, 
    -0.0448289229058683, 0.00539925845635272, 0.160623900513207, 
    0.0486003852251924, -0.0609692322473848, -0.0235145459304718, 
    0.249156799726734, 0.0892064188485706, -0.431823494369951, 
    0.144365883368402, 0.485753686894135, 0.229761756439109, 
    0.438588986460623, -0.200864882804301, -0.00322394682848198, 
    1.1826614517316, 0.555192553731978, 0.171334213602534, 
    -0.0213399422235093, 0.107823775247352, 0.278991277364806, 
    0.212090219107362, 0.100348015236616, -0.00378049365150682, 
    -0.013284761029383, -0.0451969168172139, 0.00831410333303663, 
    -0.147304391621484, -0.303600235275865, -0.0173313462535378, 
    -0.269899535915674, -0.149955627048479, -0.126432066285945, 
    -0.208235649190042, 0.0227514909165374, -0.230084283454767, 
    0.0230194367295256, -0.238023780886675, -0.0855596839067064, 
    -0.0368540821507406, 0.0321595614774659, -0.00287137805240323, 
    0.0104829547246197, -0.0361404608372489, -0.0114393779474879, 
    -7.00716525937894e-06, 0.0288295257196258, 0.0720696845031835, 
    0.0452908298637665, 0.184649414257861, 0.0280401316153323, 
    -0.0120938741336006, 0.412784537433926, 0.197637693710381, 
    0.0334841557807181, 0.179086770488192, 0.373834740043816, 
    0.0951631531673329, 0.213536025159209, 0.0942211115816014, 
    0.793762862913471, 0.162616800175045, -4.62541115856391e-05, 
    0.341452548512312, 0.490222809102626, -0.506668105610007, 
    0.616576592230177, 0.840260615863888, -0.0873746173381851, 
    -0.21710836745909, -0.0911178185443634, 0.173885729433189, 
    0.113867689543228, 0.0844424785104376, 0.0290881996133309, 
    -0.0713598989596087, 0.0482807606899291, 0.0454191860666666, 
    -0.134037616305361, -0.00661895931719403, -0.0441157573554552, 
    -0.0251290162204525, 0.00996267824743342, 0.00409673265185497, 
    0.0291249904449647, -0.0398412363639983, 0.0123967132272522, 
    -0.0048297653387627, 0.0038924953109804, -0.0166262639836356, 
    0.0380230424548389, 0.00599819593308601, 0.0161037958064812, 
    -0.0708805915102203, -0.00695047051002554, 0.0141646646782116, 
    0.00474395174929049, 0.0677938421808332, -0.038733987184707, 
    0.039575617642978, 0.0729532541801308, 0.0858200283290821, 
    0.0936539942390129, 0.0970240541790882, 0.0882146556331566, 
    0.0916588899956281, 0.110269722651874, 0.0964326500559634, 
    0.0787977982224277,
  -0.00143791184236243, 0.0869925160584065, 0.0506689012001864, 
    0.065141214528039, 0.0901471396891863, 0.0564051634540347, 
    0.0609395812280856, 0.119068537221753, 0.0995251917313655, 
    0.0283194368421584, -0.0589565126753385, 0.257030077589161, 
    0.317094248425228, 0.152431422683481, 0.000381076512119966, 
    0.24051787266507, 0.050834573073047, 0.401550562515329, 
    0.581493189473621, 0.130396373584861, 0.0178144407221392, 
    0.218628390497002, 0.715142028085026, -0.0103962640232519, 
    0.746520954956912, 0.816741994125906, -0.0318897343579421, 
    0.452516987036203, 1.02383149641899, 0.0790593556027042, 
    -0.0600233332017247, 0.00166648320270728, -0.0587320356343359, 
    -0.0136488071052528, -0.0534393555788502, -0.0357023373857643, 
    -0.0174578179919731, -0.0430009606621605, 0.0339911454241245, 
    -0.0784558617061769, 0.0509444150775728, 0.143448725949394, 
    0.111821572069383, 0.105043996734981, 0.236472192270309, 
    0.228279019408676, 0.20824969290694, 0.368103162892921, 
    0.242066297982421, -0.225282782157435, 0.438003479344831, 
    0.474542627743517, 0.0166474009833386, 0.17529760526525, 
    0.746594267491481, 0.449340386717907, 0.152344517172192, 
    0.0549008020962742, -0.359381055392227, 0.0656988036048789, 
    0.513816863734777, -0.0079808529677755, -0.194699270370115, 
    0.0768681400037532, 0.295732366440791, -0.00702257281897542, 
    -0.00527572954911691, -0.038720666950837, 0.294490810259376, 
    -0.02240102945737, -0.0624924854719394, -0.211489736095933, 
    0.0372477841609366, -0.0700875959643808, 0.0513306864020314, 
    -0.157715040399731, 0.0355543458870149, -0.0425619659396997, 
    0.0980292922152789, -0.252253031380242, 0.0650514048362457, 
    0.21244348877114, -0.105570331568971, 0.183181559845571, 
    0.351037302893733, -0.0438834719653534, 0.0268567824787598, 
    -0.122872000364392, -0.0537166752782144, 0.23771856797595, 
    0.431830702034415, 0.0793563179439064, 0.541448116722363, 
    0.761397636469585, -0.0803824243328349, -0.643718750957817, 
    -0.0763273207757517, 0.794927425480305, 0.271596666106057, 
    -0.0353047054488129, 0.170070160199601, 0.590706594790308, 
    0.137329051530677, -0.0216388687542353, -0.105992357820282, 
    0.10416340834221, 0.407696766575084, 0.345351988248461, 
    0.152376990686068, -0.0231621814525217, 0.343099394416835, 
    0.138839238789169, -0.0531406873682329, -0.127107785573113, 
    -0.106305818596372, 0.202273497492201, 0.113859001007761, 
    0.0348227861434755, -0.0787527208805498, 0.00620241152816717, 
    0.052825627997344, 0.176744322316468, 0.113309666669855, 
    0.0776312985438093, 0.141257747834749, 0.0310353788037975, 
    0.0171275065319305, 0.0627442917301431, -0.0718318295921273, 
    -0.0046523615526216, -0.0583127809595987, -0.0313695109118242, 
    0.174040486327444, -0.142472248725489, 0.0610109435004449, 
    -0.280048752619221, -0.0839846561519929, -0.109953965479199, 
    -0.0825829908682323, -0.131697717812458, -0.0116249386185484, 
    0.0664577171436978, 0.0976905016946432, 0.112048664640187, 
    0.136772444147444, 0.123003788292483, 0.130367400656138, 
    0.178725510456185, 0.137490279649868, 0.0859659598243601, 
    0.200946665852351, 0.155647578143534, 0.145378421201252, 
    0.471835398532275, 0.312362238082931, 0.0209903058348046, 
    0.0324486314665458, 0.54909384889533, 0.37993509762369, 0.21704814189754, 
    -0.201229988880111, 0.51630438187454, 0.307088609804979, 
    -0.0289507120559736, 0.397486360648036, 0.417484774903389, 
    -0.000658732569642967, 0.42337803060541, 0.559526942020107, 
    -0.033916276812436, -0.139091808362331, -0.00696840720543927, 
    0.536121259885446, -0.14633713405575, -0.136909920776056, 
    -0.0403406739169903, 0.240160141587895, 0.185312800535657, 
    0.492931919911181, 0.0483516922232809, -0.260203662580672, 
    -0.0594407946871659, -0.181907857989324, -0.107532631197611, 
    -0.151816332828322, -0.167827413809712, -0.148870507145822, 
    -0.147600764305424, -0.0840872282406789, -0.187255212874215, 
    0.0226207573545537, -0.0398323303098364, 0.0635633434248293, 
    -0.0307851820511602, 0.0445912943773527, -0.107960577165658, 
    0.0127149747266495, -0.0120591823950564, 0.0630446137462519, 
    -0.177789260352652, 0.0193626662296251, 0.0565746026000038, 
    0.0285404646823935, 0.0979093536511366, 0.145854913547177, 
    0.0768086761715359, 0.0742448095919426, 0.194964169506302, 
    0.164181391519024, 0.1599592739546, -0.118038928722357, 0.47890660433653, 
    0.281992782590972, 0.0798351933772699, -0.2011299105331, 
    0.205287948824114, 0.394836490728233, 0.419915760349055, 
    0.449000125650295, 0.248715235188148, -0.300268654824139, 
    0.487789797948136, 0.473005823601068, 0.191850494787529, 
    0.193250845331277, 0.287208045542353, -0.168603080947755, 0.164736761023, 
    0.646487390773796, 0.293912674224045, 0.382604760252394, 
    0.478805793779013, -0.11090444400943, -0.0911410194236094, 
    -0.10779608026462, -0.0207286400318902, 0.0184073154954065, 
    0.148469751988423, -0.141400086718034, 0.12442948430835, 
    -0.126598002598721, 0.234712235679783, -0.198629144935515, 
    0.138013033529738, -0.234102797933594, 0.075650248316436, 
    -0.215121721741946, 0.0288579844420858, -0.234945004606809, 
    -0.077884025549904, -0.0274665329374652, 0.0278992078997531, 
    0.00574433457435215, 0.0228809895993976, -0.0463425708787945, 
    0.00367550592850947, -0.016074236140313, -0.0264214698314618, 
    0.0868376528839317, -0.054380706797079, 0.0276934680626468, 
    0.167267741741828, 0.107693905660082, 0.013822242571753, 
    0.260804223319849, 0.246669009980633, 0.12840937615826, 
    0.0933950308479752, -0.208117149189677, 0.217018678765275, 
    0.416100448009165, 0.0528748152607918, 0.12024824603353, 
    -0.420016840137962, 0.240258590949538, 0.47117966394071, 
    0.480013816035966, 0.405056064192764, 0.112426858221724, 
    -0.301425491541546, 0.252113018932401, 0.473544556508262, 
    -0.0889965666097392, -0.167146875460688, -0.0594403800415251, 
    0.110450600137837, 0.268655522282662, 0.427178716443064, 
    -0.0262600484977962, -0.253194848630264, -0.0375197143227315, 
    -0.230791409787547, 0.0708100838089155, -0.225095242410625, 
    0.0216998112372896, -0.227180753871863, -0.075122257878937, 
    -0.18737582877713, -0.163237013091477, -0.113477802977064, 
    -0.128769275168997, -0.0138170789145907, -0.0995141326295376, 
    0.0142160220148974, -0.0900795086517064, 0.0195549095295487, 
    -0.300909861007103, -0.0708458498499223, -0.035878295557972, 
    -0.2035504688331, -0.00605168176788708, 0.0388064209906593, 
    0.0597823631889478, 0.0855274934560347, 0.100176613295893, 
    0.0857062505150723, 0.101748982216365, 0.141231080326352, 
    0.0938687051596741, 0.0441471639429229, 0.224165093992524, 
    0.171236681119971, 0.0290533277765707, 0.377691660089979, 
    0.378555566307119, 0.100923047912899, 0.0208303807795511, 
    0.506469197571856, 0.309174678464607, 0.15805680270799, 
    0.152387822817938, 0.0872465285767272, -0.171135725436708, 
    0.756969152114818, 0.265985770527774, 0.0239500489918176, 
    -0.0153242245364504, -0.245836562784188, 0.661547894182234, 
    0.332440340601054, 0.000889673060681009, 0.246536976463626, 
    0.269985651234394, 0.0974280574661649, 0.194243013456021, 
    0.319004548386765, 0.411736683057526, 0.336335509758759, 
    0.00286869865365269, -0.218792683294714, -0.00545761692829086, 
    -0.207168968211168, 0.0493356368695689, -0.312887459547188, 
    -0.0683325435703619, -0.242323028465199, -0.159468037374455, 
    -0.174035598927685, -0.0989644363875057, -0.196629064951835,
  0.285958870709606, -0.00511771079858206, 0.138939639020808, 
    0.494414321921794, 0.0836209548788678, -0.030247382298634, 
    -0.0780951835008834, 0.32551799287015, 0.255903805008354, 
    0.14863050385366, 0.154946325908663, 0.115177065907723, 
    0.0807944309016138, -0.0651272468241376, 0.0674665172253896, 
    0.652407419848937, 0.587012361472818, 0.256260967466494, 
    0.0582233704266977, 0.219438751077987, 0.580363591246082, 
    0.522941673745631, 0.293844643258107, 0.168382512004249, 
    0.197532795168482, 0.342499090957002, 0.357280782515317, 
    0.204872255226317, 0.0788737114386352, 0.414796150241817, 
    0.377728239987161, -0.0572457699077119, 0.649143395071903, 
    0.484735724631736, 0.121559452884193, 0.160629843862112, 
    -0.295080398380396, 0.0146105413859254, 0.25486423969505, 
    0.4510159487643, 0.54075303931926, 0.136608188898934, -0.106010517541889, 
    0.049491075518653, -0.23018263298786, -0.262508943891183, 
    0.426046071914677, 0.357586289852844, -0.320217293454988, 
    -0.154130272999517, -0.439740933999166, -0.0252048686061861, 
    -0.174803913642258, -0.24840647436138, 0.0810166531149493, 
    -0.216180551390395, 0.0605294761059317, -0.187026077497946, 
    0.041574154149079, -0.278110920761133, -0.0157862371512124, 
    0.0715127670667414, 0.0929430783445651, 0.15023927485335, 
    0.327537658607528, 0.274289012353496, 0.109262934525103, 
    0.0759614987862331, 0.369711699495741, 0.313994082331875, 
    0.132911435639957, 0.131214870713168, 0.517809789734555, 
    0.270508405202253, -0.026639777881484, 0.137074156865024, 
    0.568975781080227, 0.271588277863295, 0.0616810797445821, 
    0.0788399213750255, 0.337006403871443, 0.372930039307934, 
    0.250318372354166, 0.188569854019022, 0.223267242273298, 
    0.28036158991337, 0.239719339600391, 0.1206618280167, 0.0351162058961627, 
    0.418525822071009, 0.288659642460607, 0.0228319517054292, 
    -0.0303354891846935, 0.408944730213538, 0.339042120189472, 
    0.260390900814504, 0.223368477161144, -0.0990202343497222, 
    0.503531808585778, 0.281964438682405, 0.221213548051029, 
    0.300842630910538, -0.0518144980633883, 0.611045783925989, 
    0.213076761387569, -0.0863269265644697, 0.0323764534870685, 
    0.495759112092386, 0.152936382407363, 0.0294278701421835, 
    -0.0346287607993625, -0.238276979930441, 0.215615819486691, 
    -0.0466134671912543, 0.202506657732822, -0.207289021857625, 
    0.175536738370157, -0.310158887664723, 0.0574437426802157, 
    -0.250414340916449, -0.0291739674992292, 0.113857524153749, 
    0.0479406815357311, 0.054901178799452, 0.106177309384671, 
    0.12233688774898, 0.096220212769613, 0.0880113053241489, 
    0.000448997862378925, 0.0174584343715814, 0.066513079105587, 
    0.113233726762879, 0.122619777069282, 0.142673551911543, 
    0.139231420712436, 0.0542024678798972, 0.191218376449866, 
    0.278664866779135, 0.0294223075515361, 0.157448617454706, 
    0.48319802933482, -0.066217190474987, 0.331134796143532, 
    0.589971671293716, 0.166023009433501, -0.307217476524185, 
    0.278474592702962, 0.51212592092884, 0.287785686608327, 
    0.236705374065543, 0.206410600029345, 0.347996085869848, 
    0.270230087935367, 0.0292460869156871, -0.0571031671090107, 
    0.0757963315400486, -0.215504955028391, 0.0284514615915274, 
    0.0397775989534491, -0.300481814535724, -0.331379103262994, 
    -0.214574704038273, -0.0256050059679412, -0.321492296032637, 
    0.293741275043775, -0.196112335955196, 0.0839346255922571, 
    -0.318278810202731, -0.0513112516746456, -0.29452434363367, 
    -0.149288646524628, 0.0577314274511123, 0.116754025414267, 
    0.0721178622996493, 0.113941682306699, 0.0761380509140977, 
    0.11153539356271, 0.112070047750435, 0.0409911016483501, 
    0.0792058258812716, 0.091777348834161, 0.0934057043245535, 
    0.0974943807429955, 0.0963424969511079, 0.101357967471559, 
    0.0908390038636969, 0.0820713948992217, 0.153880316357583, 
    0.141186432256376, -0.0763413414057668, 0.225003424573946, 
    0.328003781150785, 0.152319198467413, 0.0487477643780203, 
    -0.0204199533732813, 0.101492919913477, 0.520926843688557, 
    0.31785103623529, 0.0752072571861441, 0.157127971244373, 
    0.391970733248296, -0.282585002099257, 0.377984148689357, 
    0.462165992267746, 0.758962094938995, 0.517444264483901, 
    -0.172796256940538, 0.532845728520719, 0.573498522508288, 
    0.152289289938801, 0.124897768453599, 0.585021420832064, 
    0.253137828623059, 0.117044965624492, 0.030223751098744, 
    0.549897546338971, 0.169080857878294, 0.0748313658743671, 
    0.00612769170575045, 0.474479336881495, 0.143904442006155, 
    0.10204618195422, 0.0696853139324993, -0.045915317774369, 
    -0.119312850451634, 0.239285881451639, 0.0493791467797555, 
    -0.0720746731104514, 0.0986775513156059, 0.193163424881244, 
    0.0730825784685848, 0.110593406760215, -0.0640492953781658, 
    0.25655563303169, 0.264990319280702, 0.0813296329308794, 
    -0.0154535961110822, -0.0136099339874394, 0.509869639639572, 
    -0.0362323434757304, -0.0765127833297894, 0.0246760970312744, 
    -0.0474605213700152, 0.0286420237218925, -0.0328266462403129, 
    0.0188146960488608, -0.110727290938726, -0.0239878334373988, 
    -0.0292080128623361, -0.0950951874936681, 0.0267229336846519, 
    0.0795424278133733, 0.0814710701970004, 0.0838777671469129, 
    0.109013983564984, 0.0904539433132498, 0.0628002421428625, 
    0.190386184061002, 0.063922571044009, 0.0216583517112995, 
    -0.288832466599352, 0.271809453751612, 0.403302758498568, 
    0.398371298159443, 0.247025759428044, -0.2388213707069, 
    0.140748979018932, 0.467325767707418, 0.476606627672361, 
    0.283010035473103, -0.371508248756077, 0.314709889465525, 
    0.50924257586056, 0.0366279095430287, 0.17351103876639, 
    -0.00016611252866694, -0.459023698568423, 0.299759636649156, 
    0.424583136219014, -0.177679065664878, -0.126626401177356, 
    -0.136251597030073, -0.107359873244229, -0.142030118028488, 
    -0.109384481227018, -0.116248596349947, -0.0457212534624379, 
    -0.103144711058022, 0.0864835297327578, -0.210749755857001, 
    -0.0121053930937293, 0.318972214973153, 0.136751320830946, 
    -0.120042851682669, 0.0201554024219661, 0.484410475274899, 
    0.22807471860077, 0.0699459817327259, -0.0884045378491149, 
    0.150806570622335, 0.388383848071033, 0.322039041377729, 
    0.16273261256667, 0.000412949773589577, 0.234985885224852, 
    0.437200689930151, 0.187232426207467, -0.00760112836054075, 
    0.331411525696334, 0.361783989252343, 0.0908101249096635, 
    0.0427101708958964, 0.019156670627132, 0.0364679400813369, 
    0.0281108356476239, 0.0319063630469491, 0.00855503006477676, 
    0.0291220516554192, 0.0395852903993808, -0.0275767034802873, 
    0.046950499918761, 0.148989864918137, 0.147590322476757, 
    0.0680374003355078, 0.123719248463643, 0.286884652358885, 
    0.151959522239498, 0.0107066595747543, 0.274831321685123, 
    0.359626973274253, -0.417595763137548, 0.156997380354734, 
    0.85536517383565, -0.0547714949420064, -0.0391183812332618, 
    -0.0873773179296716, 0.381863026360934, 0.0798208562097376, 
    0.917202632473684, 0.507707715668495, -0.219180963200625, 
    -0.108202893500161, -0.0901457953686237, -0.0795025470120569, 
    -0.0155813112775975, -0.129702489784788, 0.0482005216903352, 
    -0.0125391593539707, -0.0281293096513547, -0.0266110392258162, 
    -0.105904007906828, -0.0585920973352603, -0.217032094201813, 
    -0.0614367796985714, -0.25794001449238, -0.203548910806421, 
    0.0567330511930079, -0.0640491506860716, 0.152148996948906, 
    0.0355978491540687,
  -0.0269585577060965, -0.115745863104457, 0.0755184724482692, 
    -0.0924265261435171, 0.0569973816156752, -0.188931122979749, 
    0.0240609393273247, -0.131796935881371, -0.00753312690012117, 
    -0.178845033029134, -0.0528123722033693, 0.0167309287017387, 
    0.0117226068942932, 0.0218023011421503, 0.00483352882025297, 
    -0.0234859785198558, 0.0243877031969805, 0.195305104341226, 
    0.0581562116611532, -0.470041605532428, 0.16927401377616, 
    0.459360156706025, -0.0488836034035929, -0.221250030128606, 
    0.193963274047873, 0.587587233553956, 0.11102015137373, 
    0.971152068870976, 1.05838420191876, 0.0802677278731947, 
    -0.0907501049202414, -0.0720755367674328, -0.00650801092348335, 
    0.158030333890115, 0.157403869682008, -0.0611773334980028, 
    0.193385179668551, -0.10354898761712, 0.0587993241120102, 
    -0.100493892111777, -0.0158980658671507, 0.102225672990805, 
    0.182376682486006, 0.204050807945185, 0.181351252691718, 
    0.18915625118658, 0.281118295138224, 0.275925664998321, 
    0.218349135609151, 0.205458586408622, 0.146283183448947, 
    0.128093793350188, 0.121422912282998, 0.112054568039694, 
    0.122846132255873, 0.127945327103625, 0.125197702299249, 
    0.136505549616113, 0.130376854759276, 0.0866023710346401, 
    0.0671566148540037, 0.203215860328402, 0.218669208304506, 
    0.0722322118700257, 0.0930401714243773, 0.35036828093654, 
    0.303464275269021, 0.26614345500375, 0.279677970208084, 
    -0.197976570579719, 0.668668877752797, 0.326627909848243, 
    0.0442864141300862, -0.0313269761943414, -0.390124055362145, 
    0.0959354556290129, 0.723605310744167, 0.513701649388933, 
    0.163331317163027, 0.00952013732070086, -0.253507615041579, 
    0.346247514923132, 0.41424905120876, 0.240420629890487, 
    0.0075684830541624, 0.559633360159916, 0.0774749950029098, 
    -0.208815725517884, 0.134515136315509, 0.433858658384989, 
    0.0265600150845379, 0.0182291249478671, -0.0380035303494901, 
    -0.0665366536348609, 0.0990195459374697, 0.354603560464816, 
    0.272529656817463, 0.0759908535177826, -0.238101897018456, 
    0.0340133487016602, 0.370529914056694, 0.192150060583027, 
    0.0981005638351542, 0.681566380125371, 0.0885303615054355, 
    -0.0139896775752707, 0.117764942283871, -0.0902468279468821, 
    0.378269929148804, 0.615618000352326, -0.011983097826273, 
    -0.081056664145982, -0.0685338091040128, 0.0223635914706273, 
    -0.100306676167694, 0.0222850396410973, -0.121489981696768, 
    -0.0635888731120556, -0.108129035023571, -0.0594712581440152, 
    -0.1654272140928, -0.158545561353571, 0.113748223116114, 
    -0.117700335885399, 0.0491971188529976, -0.0351066065243732, 
    0.0434839408767293, -0.049296421658677, 0.0633308509459369, 
    -0.0765332424640904, 0.0866384920228248, 0.0204804910656918, 
    0.0391293379279105, 0.0260698629070316, 0.0375023413356958, 
    0.0228825014387854, 0.0319760266202701, 0.0418355698616104, 
    0.0488554599419411, -0.013776934056579, 0.0743463667094252, 
    0.104996108016913, 0.0908638899194295, 0.158450614371759, 
    0.196734152220598, 0.0862742020381325, 0.156985334881477, 
    0.357634372586084, -0.0867236584585917, -0.188989917096659, 
    -0.105398052033501, 0.525365971939771, 0.116278861759139, 
    -0.222321419022691, 0.137810952661036, 0.522339184643706, 
    0.463829318424977, 0.278420459403182, 0.121410378186392, 
    0.011122762917033, 0.512944680395344, 0.208237712301684, 
    -0.247587548080357, 0.23740987053773, 0.623837872314704, 
    0.209839208307369, 0.164793428247552, 0.366790061320692, 
    -0.170482803360683, -0.260804131730411, -0.310350595212749, 
    -0.181842931354504, -0.23079280482525, -0.389163026057443, 
    0.140627785494963, -0.093275586267001, 0.139803426642173, 
    -0.08716138192061, 0.0899927609964452, -0.339409934890912, 
    0.0166344487310647, 0.019496696767819, 0.152728169427326, 
    0.214361256137906, 0.0923783922841808, -0.0122224789927237, 
    0.376926641805679, 0.304541955899546, -0.0275653551016742, 
    -0.0291654516446684, -0.326153310544915, 0.153093979988297, 
    0.579411711143573, 0.322852133885423, 0.135817624010288, 
    0.302874278622033, 0.457920635536914, -0.255341437277567, 
    0.747433713195452, 0.501169387587709, -0.0656284331465017, 
    0.03733961448535, -0.252441593352359, -0.0564664296849718, 
    0.571819462979149, 0.148548208983713, -0.0516176593462639, 
    -0.0784287219066311, 0.53167085760235, 0.175922940277573, 
    -0.0970095739858781, 0.126091953436631, 0.317204381391324, 
    0.131677589152882, 0.0902913555935433, -0.0686591946448263, 
    0.350550988640173, 0.169820262208281, 0.151263367951852, 
    0.20201648664499, -0.226396769577204, 0.390390796376666, 
    0.273814981453073, -0.0296926464692108, 0.30242932456795, 
    0.357842604303955, 0.01289419442735, 0.139838837338572, 
    0.529466632377008, 0.185158211214639, 0.0359637665774885, 
    0.0705530710351819, -0.0804065440023971, 0.11098300520355, 
    -0.0215826452591641, 0.125999603818795, 0.331395360715563, 
    0.0198660585659795, -0.00978595513002678, 0.00754821851907277, 
    -0.037937996482757, -0.16211381294419, 0.0585754912526254, 
    -0.0517295733032892, 0.0643049493042831, -0.0649216455604841, 
    0.0910723491930399, -0.100527785998102, 0.0977310040609072, 
    -0.131252824446444, 0.100343012234888, 0.0264205369269362, 
    0.0480484720137436, 0.0210469118672095, 0.0343314791152471, 
    0.0337602027063555, 0.0543101497589444, 0.050898281619551, 
    0.0798220279097055, -0.00546684036073639, 0.117918012625128, 
    0.122646470114197, 0.0511072433900743, 0.063393556059973, 
    0.358792447084981, 0.124753352159787, -0.281658905357609, 
    0.170264449120165, 0.502688504987184, -0.180577727817472, 
    0.217153215065422, 0.796581948417368, 0.0858847225489421, 
    -0.44736496731545, 0.316386626974542, 0.682631791552817, 
    -0.00387003414301336, -0.0316194531754175, -0.0617965729681412, 
    0.239418710456198, -0.129996561495413, 0.275901969218875, 
    0.782972322857089, 0.24605532185799, -0.044263725997041, 
    -0.118939716037522, 0.0220130563574668, 0.560928146670064, 
    -0.185241522585577, -0.0416725477589749, -0.116792641867484, 
    -0.282513258978035, 0.152353309637014, -0.257064842596945, 
    0.126801520978995, -0.254437324824363, 0.102546167003318, 
    -0.300495187467598, 0.0312955199672643, -0.272894609522807, 
    -0.0473805599923488, -0.0217676438413853, 0.172923940832798, 
    0.114569205361249, 0.027024636056666, 0.181767309763826, 
    0.140050866892784, 0.0452888895497694, 0.221907491724323, 
    0.123108105727098, 0.398238366688874, 0.423541621675694, 
    -0.367468854374347, 0.528443047370612, 0.565068213980236, 
    0.132426488032521, -0.172996185657454, 0.679200931609322, 
    0.514535478771565, 0.208496803044184, -0.156999525412907, 
    0.561032453346925, 0.283601260259436, 0.0410448902178551, 
    -0.130121312479465, 0.315882495625499, 0.524063642742854, 
    0.181628248601245, -0.0432715488179025, 0.173830065204832, 
    0.186010127294811, 0.0778128515683639, 0.16257981484999, 
    0.250777596506595, 0.110066540572523, 0.0293878487399884, 
    -0.0302563234339836, 0.217549406305486, 0.0538815412576061, 
    -0.225102260744746, -0.067549764645883, 0.443560166521665, 
    0.241517189963679, 0.156259658081423, 0.16366116233714, 
    -0.167094409978203, 0.17687396544718, 0.262405961153324, 
    0.465343190587196, 0.501175311533914, 0.0754013251059635, 
    -0.0229445711370049, 0.0210753795770922, -0.0199179970022339, 
    0.17517486094773, -0.00442673068319174, -0.057309467071821, 
    0.0629003755615914, 0.0892216331380065, -0.00245392278851224,
  -0.0308315160518606, 0.110718644357766, -0.116295073162941, 
    0.0901609517429317, -0.0868655093536579, 0.0677181017479429, 
    -0.332767286431523, -0.00495332268680446, -0.291157487909227, 
    -0.221764338818846, 0.0162356745608639, 0.0599224765924255, 
    0.118390266028409, 0.214415217463067, 0.250282292949461, 
    0.227926565602445, 0.208235781246631, 0.214201347402611, 
    0.243500073946294, 0.280767681647195, 0.313276342025374, 
    0.301127074233776, 0.282326482553791, 0.273265410691655, 
    0.258343402376637, 0.245466124366033, 0.266968928051094, 
    0.270047356918679, 0.236325009052204, 0.296944431192909, 
    0.357203833162182, 0.20735764398416, 0.0326843666567506, 
    0.241112373219013, 0.352023109761003, 0.0968026081911457, 
    0.175750912591907, 0.509350924978962, 0.259147496348302, 
    0.133463466231368, -0.0117018070347645, 0.537899977575409, 
    0.337418088146706, 0.114092377905407, -0.198106831874027, 
    -0.0591069843820856, 0.407123931901805, 0.348809539016261, 
    0.315597358097847, 0.26630574599012, -0.0116649602578423, 
    -0.188541157188564, 0.200332509362635, 0.365489105628434, 
    0.0963569198104868, -0.186991705986971, 0.244995935636216, 
    0.205510651969571, 0.0585079541062751, 0.00457543745436234, 
    -0.0766147405578396, -0.222942705720949, 0.0464079340315275, 
    -0.0915230630289738, 0.0385014775594392, -0.223103650186257, 
    0.0425432722868304, -0.179166584388716, 0.0198081699452113, 
    -0.292964098290477, -0.0416946029513125, 0.0333772200609847, 
    0.102435573569448, 0.12637324255459, 0.125042904066525, 
    0.103193036815957, 0.111626435965745, 0.147786347679802, 
    0.113373361126264, 0.0729134680343191, 0.201526408769455, 
    0.171282119538278, 0.0876202049776675, 0.305009991549545, 
    0.333654292226855, 0.0989658218418805, 0.164718534333851, 
    0.540895036078272, 0.132077552346134, 0.00985743318574582, 
    -0.199387081433291, 0.0246261441655832, 0.639252531384125, 
    0.196001440469149, -0.0679632498104842, 0.0802747480859371, 
    0.273539620311049, 0.197343104028133, 0.632452439248229, 
    0.415271690804323, -0.0798491498030045, -0.296579069055949, 
    -0.026710008768316, 0.533342159872075, 0.162822088703965, 
    0.0870867733073395, -0.209676566134273, 0.28472546742075, 
    0.0123451159193943, -0.223986836872047, -0.307254770281511, 
    -0.00847854550848144, -0.246703590566811, -0.0123382360664276, 
    -0.260513950164772, -0.0443241227196413, -0.237758454194045, 
    -0.0856094253933771, -0.231807518280478, -0.158411577152105, 
    0.0410885506789825, -0.0922540163590575, 0.0855800837185151, 
    0.0020820167208369, 0.054229651789137, -0.0249079797019929, 
    0.0267544435978726, -0.000847465245170889, 0.0603298419914956, 
    -0.103001192764234, 0.0343910518506946, 0.0809337699869455, 
    0.0600395650323978, 0.0886447155497834, 0.130954425305791, 
    0.166496969986317, 0.213486789046932, 0.104352071161457, 
    0.0119096451255254, -0.133245929202625, 0.566813916908297, 
    0.151795586729469, 0.0013932555477669, -0.188942904515136, 
    0.00106918699139429, 0.71836607503726, 0.208554705909477, 
    -0.120670252043839, 0.0958879509518793, 0.540529145795784, 
    0.195796933290501, 0.0823774911501601, 0.325320495134333, 
    0.123203630874631, -0.0539255974974269, -0.150901028029196, 
    0.300696053467971, 0.738156408680634, 0.101845637869708, 
    -0.145585682961468, -0.08616213818536, -0.214441742365018, 
    0.0610391550223162, -0.229801157908622, -0.0609515482707558, 
    -0.213342960793281, -0.14209798350219, -0.0156483614508569, 
    -0.17102910109101, 0.108087054570785, -0.168150907634031, 
    0.0500208425431205, -0.132982483079688, -0.0366169591938871, 
    -0.111212441924642, -0.0620123001365817, -0.131382243639123, 
    -0.0852017324001694, 0.048782622031843, -0.185854911247813, 
    -0.0331774843909312, 0.113105020766652, 0.0528001931283005, 
    -0.0133326164194232, 0.141897472764843, 0.14303092316095, 
    0.0194410192575424, 0.200009486279703, 0.278273075762187, 
    0.0467706336218363, 0.121818339840287, -0.182215409248453, 
    -0.201063556826775, 0.638498619567835, 0.390984005376723, 
    0.158897015873208, -0.24942508588439, 0.235704500550794, 
    0.283582804867505, 0.573035667122769, 0.494644155456206, 
    0.161778116674812, 0.7749399507335, 0.681027214223244, 0.328634587710373, 
    0.0893948626279887, -0.358943631074552, -0.201090148314563, 
    0.752774938681779, 0.0843936960970425, -0.188908798948843, 
    -0.0482306701433765, -0.0638543655724524, -0.217771490067817, 
    -0.240198569525378, -0.168819671503594, -0.304464102606823, 
    -0.221578151129251, -0.109531178609652, -0.271732004256059, 
    -0.108222973773665, 0.0232690501490619, -0.0795638866091316, 
    0.0179306349462166, -0.0984796679209184, -0.00290537421233832, 
    -0.0930261126188105, -0.0427923922662844, 0.062662740260137, 
    -0.132718902422374, -0.126893350130949, 0.324802035611421, 
    0.22783592422254, 0.0417667303083886, -0.117154326269745, 
    -0.0936644970280019, 0.457586082164509, 0.240998843462898, 
    -0.0136490050278515, 0.271513841198669, 0.404215522649551, 
    0.201707740025118, 0.0813664298218316, -0.041958082444032, 
    0.228425725316134, 0.290712233304759, 0.108743406035444, 
    0.104080441421112, 0.389806224182876, 0.168520378733889, 
    -0.0292415233933438, 0.00594369948811047, -0.0780512873297208, 
    0.00985127117604591, -0.101424586053103, -0.0311646916973072, 
    -0.174993572841301, -0.0866164764419849, 0.0558831178235553, 
    -0.185566926895198, -0.025935600346831, 0.190070079488104, 
    0.062280717545506, -0.0401013287154459, 0.00711265390188036, 
    0.338137211746628, 0.166565414962238, 0.00942572496600094, 
    -0.0297830135034559, -0.0856747841980332, 0.852186101211963, 
    0.169672600085456, 0.195163118642953, -0.448768821346603, 
    0.168519505456698, 0.75276703173244, 0.141789064161919, 
    -0.338806652109031, 0.416457540251208, 0.239819031968603, 
    -0.445588614209053, -0.176987613487653, -0.000806313973890221, 
    0.372187155739676, -0.167633853933693, 0.0411064539150439, 
    -0.0735646224289139, 0.261103886745403, -0.171251224384814, 
    -0.495320276851777, -0.069803349143619, -0.342817672488811, 
    -0.11040271851943, -0.208449164466599, -0.242344697271235, 
    0.012861663564671, -0.241961290132019, 0.0298794187143596, 
    -0.401565863816128, -0.0530868367030335, -0.07549061888139, 
    0.0784900121357163, -0.141627867609356, -0.0399766931367201, 
    -0.00164136045692792, -0.0779875886851989, 0.0277986737611595, 
    -0.0342560596084068, -0.00100031466717043, -0.0199354913864658, 
    -0.0907801022192546, 0.134392587387392, 0.207580860230775, 
    0.0310445366649491, 0.0208514339848802, 0.370245212821854, 
    0.218763876351417, 0.0794072123421648, -0.0919256064663506, 
    0.362349370137607, 0.316223309722706, -0.159858794145464, 
    0.264805346427567, 0.592687246422728, 0.206310955447864, 
    0.128628869913662, -0.250012938419045, 0.173375340278312, 
    0.441786038754179, 0.216882917717252, 0.162030002792865, 
    0.446516028981216, 0.248661424465538, -0.0722170354644954, 
    0.2407469261066, 0.604203562734209, 0.278520405449622, 
    0.0891007846123879, -0.14129132494056, 0.178641866766811, 
    0.493692771500739, 0.38533451777583, 0.0967352522136208, 
    -0.181510649086963, -0.138110399230176, 0.391803274504637, 
    0.403629812592988, 0.163299268069398, -0.154960759283276, 
    0.145179018993111, 0.295509998794927, 0.203359799653708, 
    0.236676782647963, 0.0791775978114613, -0.118441468585967, 
    -0.150795981238033, 0.287360987461603, 0.140807087943729, 
    0.251988592252639, 0.256264545916288,
  -0.192877979155758, 0.129792671263589, 0.468866142932346, 
    0.157289399881864, -0.0350503189790081, 0.0481816640859144, 
    0.391349874178212, 0.134401416248516, -0.144507527712077, 
    0.144746256996518, 0.895894440008734, 0.188459448367463, 
    -0.122947697236746, -0.0892907011221983, 0.6979095092196, 
    0.283039990092238, -0.164032666235804, 0.597410934001866, 
    0.961265065711329, 0.449770088713819, 0.171596435617997, 
    0.283708920624618, 0.276194111994093, 0.158442430004571, 
    0.18526227277881, 0.319946624217571, 0.264270698546028, 0.13463855154696, 
    0.0686321272506175, -0.0859544824998985, 0.454380424949603, 
    0.18008714692143, -0.00909439050204366, 0.00277427554706892, 
    0.470870044896225, 0.13073049383593, -0.132749743691861, 
    0.19899333327289, 0.284543990554048, 0.0494497454187409, 
    0.402185368438474, 0.470421253692063, 0.127548043968502, 
    -0.0322685529701469, 0.238486479522327, 0.185844252073504, 
    0.317260108782403, 0.433796269441395, 0.257131367478, 0.0735094367018483, 
    -0.243424085775257, 0.0780200804642867, -0.204949844765001, 
    -0.0287514819799446, -0.366469914460192, -0.204473424420256, 
    0.138103437468608, -0.237714105587408, 0.173778172534936, 
    -0.110981444101764, 0.14999761784398, 0.0533039061929251, 
    0.0524430505345818, 0.0897937133967783, 0.0905007707367518, 
    0.0265737465184717, 0.0655504178734443, 0.101376358649194, 
    0.0825660712440665, -0.00150829421223232, 0.0543586921153504, 
    0.128376732114945, 0.143056094548163, 0.130740107661182, 
    0.143549338572978, 0.193298177557296, 0.26461581483059, 
    0.156053244919038, -0.0884644031300839, 0.135906810070393, 
    0.489121400870145, 0.15786867944998, 0.14169430139779, 0.767870980581853, 
    0.228729365643813, 0.0115070063391169, -0.0286930093281374, 
    0.610709360188246, 0.351025429977933, 0.17443591150531, 
    0.222665674101363, -0.477670000058398, 0.52414724104043, 
    0.255295622140138, 0.0352277015879964, 0.693970319130206, 
    0.116346992569439, -0.348261403217088, 0.274861649094432, 
    0.339258449870097, -0.350509579093931, -0.109219332679656, 
    -0.281239172125558, -0.142457173255832, -0.125719917884217, 
    -0.126622842470667, -0.191195490393516, -0.0957572560166086, 
    -0.329765102107225, -0.0747063442238619, 0.0570826127106361, 
    0.0823990758880568, -0.302342389727867, -0.00953616292610529, 
    -0.0672185155061205, -0.215826951719394, 0.121604723890049, 
    -0.0387242273103916, 0.0778823423847408, -0.225630560829853, 
    0.00270553206387873, -0.0105619391926157, 0.0672949273115298, 
    0.11489622033511, 0.059976650807067, -0.0115877919578799, 
    0.178992989653328, 0.117346423339321, -0.0210688803511814, 
    -0.00427582863511296, 0.22917216068391, -0.0517621871544721, 
    -0.172121009649265, -0.0626343497046817, 0.667336835388889, 
    0.382210223943432, 0.0620777559724555, 0.587551473828622, 
    0.537722405018593, 0.347457297121594, 0.264012571997578, 
    -0.135621809315441, 0.603636501182098, 0.272771435830223, 
    0.0749523540294269, -0.201860753745313, -0.0252077137871517, 
    0.516675085755694, 0.344825246960259, 0.167070770508324, 
    0.192440659064072, 0.153831398659576, -0.151879131348293, 
    -0.127821752289468, -0.0385480702599513, 0.0480091711695679, 
    -0.0390821953697098, 0.0120967372202713, 0.118756727772419, 
    -0.154031648250357, -0.0171459185376235, -0.0983653865068663, 
    -0.00689160372387737, -0.0616152417872212, -0.0461539660139168, 
    -0.0633935149375717, -0.0623194018964804, -0.0672788262697957, 
    -0.0267016824854033, -0.0304885679681599, 0.00224591313882121, 
    -0.0421941042971233, 0.0775351522214777, -0.0861166994106518, 
    0.0554327732212315, -0.123934969816819, 0.0207543711291906, 
    -0.15341983912841, -0.0348951255892013, -0.159755269006975, 
    -0.074447200911033, 0.0206825878228177, 0.128348601537322, 
    0.100109455075297, 0.0563084342531933, -0.00564638273021864, 
    0.0803891345711786, 0.233212470750427, 0.105622951687964, 
    0.00415874948389571, 0.623014644824079, 0.148203713506094, 
    -0.0561659346776481, 0.148442196135347, 0.692615207768105, 
    -0.204573944832772, -0.0310085739430413, -0.295507485677578, 
    0.287702430096904, 0.542928710955907, 0.298846425929701, 
    -0.0538119124391686, 0.521529507319324, 0.217059405208852, 
    -0.0402566239868607, 0.0227631376454735, 0.539081117488958, 
    0.221587523621349, -0.0404990479071118, 0.464142446694056, 
    0.292940502752337, 0.0638755603183783, 0.000347018955541428, 
    -0.0616258314182447, -0.0571111986569044, 0.104229189554483, 
    0.0456424352790781, 0.39070369032235, 0.085481080526359, 
    -0.112932194217495, -0.0818812223621661, -0.116048408386693, 
    -0.0549090346169095, -0.0688942080770569, -0.0841422304278192, 
    -0.0722366488127595, -0.0731525580406329, -0.0267369160962624, 
    -0.0787133459509458, -0.0148351510286456, -0.0400051865854493, 
    0.0508464486270306, -0.0655624632399367, -0.0081204551223089, 
    -0.0422374370080424, -0.062494610570822, 0.0810194507639941, 
    -0.0157450553127656, 0.0875990689939098, -0.0860474945023182, 
    0.176912050333738, 0.171081040688172, 0.0446592809498118, 
    0.0617369459572228, 0.211745446936612, 0.277325687625175, 
    0.163842644332074, -0.103711586472405, 0.320846939728329, 
    0.36964831177041, 0.222729679612898, 0.0316049600922539, 
    -0.253672414825889, -0.327295318742832, 0.742229758935182, 
    0.369514467085392, 0.0479019394156675, 0.702811405488532, 
    0.320960060628919, -0.384977653573181, -0.250736305278133, 
    -0.0658571971651706, 0.0732318687283765, -0.078418492561914, 
    -0.068642829398788, 0.0219190786142626, -0.127030781154496, 
    0.00548380533922625, -0.107479126189282, -0.187317050035717, 
    0.0150331264861994, -0.107855273651622, 0.0258004761000363, 
    -0.127534687824756, -0.000590010516222206, -0.0991243866394086, 
    0.00459014178208883, -0.11799014582809, 0.0480128904424331, 
    -0.0976538707585295, 0.0481826703788755, 0.0180264852347706, 
    0.0464834431695929, 0.0246181692750961, 0.0400791488799657, 
    0.0217526954547705, 0.00642083410999446, 0.0861562725986655, 
    0.0757162181503148, -0.0495485339573154, 0.0400708943848831, 
    0.2168151898963, 0.151099450625332, 0.057007043011133, 0.185405214262219, 
    0.35886575097734, 0.21770641565818, 0.0775012254029228, 
    0.0867818049310516, 0.445844513877229, 0.48370119467332, 
    0.296006043270821, 1.03916694676439, 0.216277307474228, 
    -0.140142313911395, 0.41496602574956, 0.535770732010048, 
    -0.105750710794174, 0.93579493381814, 0.727351901039409, 
    0.0705702446489144, 0.0254443295572102, 0.0611457510629173, 
    0.138193641564092, 0.135037945701882, 0.0733606328110797, 
    0.0907125540025292, 0.104685986777419, 0.106971330196879, 
    0.0684304163169464, 0.223543880897287, 0.136277966734231, 
    -0.0364719667285004, 0.444671700191943, 0.241933437339678, 
    -0.0160685342411337, 0.210143329956274, 0.307185849917027, 
    0.158036132256756, 0.49421128048833, 0.296616616665578, 
    -0.0260400870077356, 0.0612666550177313, 0.970005552206631, 
    -0.279129571305429, -0.0130472657883401, -0.383741539313836, 
    0.336575966151268, 0.610127723390132, 0.263947815022527, 
    0.0184825436265427, 0.440179344731886, 0.143009167287359, 
    -0.0452959408714012, 0.217971558391233, 0.206806939047106, 
    0.055693173988366, 0.07751272739536, -6.02247751858298e-05, 
    0.198281826660585, 0.0834004519394237, 0.039042445194511, 
    0.0319846496958021, 0.0315345953866838, 0.0374386494444786, 
    0.0386426045616579, -0.0213315991846428, 0.138728758523822, 
    0.048493936274655, -0.0817818388901166,
  -0.188992413697223, 0.0220539113885197, -0.220272390674407, 
    -0.0640580415307227, -0.167727502720517, -0.129624086601296, 
    -0.233945132657379, -0.0863201181502067, -0.21385283764771, 
    -0.00210348493254189, -0.146513941466558, 0.00620618466748805, 
    -0.0993056056384362, 0.00445643064587216, -0.147267744362254, 
    -0.0645600287416828, -0.0701898966486585, -0.183825314907037, 
    0.055164180100223, 0.0435743593890144, 0.30927910041467, 
    0.0494657885591622, -0.0910350908271453, 0.37629151639406, 
    0.292044868058375, 0.120241846979045, 0.0154274489676095, 
    0.44981938913128, 0.108088212151745, -0.489837589434066, 
    -0.0231303629616993, 0.719251610131878, 0.278830438707369, 
    0.177436272534285, -0.378267898408676, 0.114193830269625, 
    0.664615245991901, 0.187850579763167, 0.0861351165307639, 
    -0.240323389323731, 0.542083642879502, 0.32829691472796, 
    0.0665909683313343, -0.221659079243603, -0.10946310871895, 
    0.57668403781236, 0.220179167849571, 0.122224073036545, 
    -0.0813437037062502, 0.597444743855044, 0.142409456816573, 
    -0.0323533336303475, -0.0344841785950218, -0.173183194825546, 
    0.534305726266789, 0.150452767375176, 0.25679881224529, 
    -0.369916104508148, 0.172209155162612, 0.311106478058428, 
    0.17525891935312, 0.166492444045786, 0.0309238055337403, 
    -0.0241857734984745, 0.246221348726684, -0.00929111382463237, 
    -0.169132222278221, 0.0965230193574945, 0.10995409666588, 
    -0.149074223190701, -0.0578295557448558, -0.073517313545922, 
    -0.0213750762077648, -0.0912872648973812, 0.0384505384417062, 
    -0.107078570387475, -0.0202905422675393, -0.0683228149151996, 
    0.00304756276724191, -0.0773614793363538, 0.0139582117364827, 
    0.0758153999499357, 0.0983159956489149, 0.105309061584066, 
    0.097318188123248, 0.0677087564484276, 0.0740600064658085, 
    0.278382659668996, 0.128893103553341, -0.219935375737643, 
    -0.0322063956573339, 0.436246538239134, 0.353723580012567, 
    0.182916874108971, 0.0710469821026795, -0.234722099855843, 
    -0.0698181597354223, 0.463366939826755, 0.633398939210941, 
    0.248159291549715, -0.19217729524855, 0.250626593236503, 
    0.481986175218243, 0.143826328559897, 0.00918898754671441, 
    0.642419461110061, 0.605236515548147, 0.224924737663178, 
    -0.213687952583918, 0.149429437353323, 0.545407108761006, 
    0.118329361557912, -0.0533411016119832, -0.0877944360213376, 
    0.0467400447650883, 0.462785393862329, 0.437589922565361, 
    0.173468788465748, -0.267559126352747, 0.363481786623199, 
    0.498674285517276, 0.200053350788991, -0.028459204584757, 
    0.487002954707745, -0.106033576818748, -0.242658196886452, 
    -0.192892937401368, 0.140844278310597, 0.298569894336579, 
    0.336474580640719, 0.149044322680082, 0.15996270700482, 
    -0.196428989056035, 0.205097990139044, -0.335946659367945, 
    0.0600023320052598, -0.357252713638742, -0.100223558783167, 
    -0.195899346610724, -0.192152655162728, -0.0332878202448519, 
    0.092312283892422, 0.0836787215574143, 0.0963013663309515, 
    0.100433499993222, 0.0795824465884414, 0.0503182357553677, 
    0.0896326454617672, 0.103529780838223, 0.197974678613291, 
    0.261337858977274, 0.040124545786838, -0.12161435389118, 
    0.15464539707961, 0.411728683457295, 0.499504339638611, 
    0.260398064067891, -0.0302196474548129, 0.264122365888659, 
    0.384389631283384, 0.0397187742813512, -0.169421287308935, 
    0.263222730095949, 0.996180208847323, 0.13864726709596, 
    -0.158236723839216, -0.22571084028285, 1.11196733719304, 
    0.0655987514967139, -0.0436554227528975, -0.152896631645449, 
    -0.233474409853003, 0.0127831886183018, -0.232104296536985, 
    0.0110128410664111, -0.185296370105989, 0.044320305007877, 
    -0.150898364972809, 0.0631526240504062, -0.210229173317562, 
    -0.0115828841216268, 0.0937711334826016, 0.15218533719183, 
    0.181228631677596, 0.19327576049583, 0.184336027219144, 
    0.195088417520931, 0.224541795095035, 0.165299269048776, 
    0.0767206009277546, 0.286418536506347, 0.39229690425214, 
    0.193205928506644, -0.0494523396930187, 0.200072683608023, 
    0.566369670290489, 0.27410455158956, 0.0841107823947871, 
    0.0317452141476929, -0.0954124134560805, 0.303462620498983, 
    0.67503868190453, 0.31032750431781, 0.0629448593831147, 0.67592389614193, 
    0.265512672274151, -0.439913084805211, 0.198754416112853, 
    0.731264464309864, 0.115520305184742, -0.0652527545458423, 
    0.00163597736114904, 0.0264404503483569, -0.105872530018484, 
    0.17732901607735, -0.182658456158137, 0.146795411344258, 
    0.193234743529584, 0.0342974025341549, 0.0196087365127612, 
    -0.0410722094023677, 0.0457979560953133, -0.0889557448737515, 
    -0.0122756235600305, -0.0531635616871454, -0.0648528404986922, 
    -0.0198383855000074, 0.0867291873961349, 0.124903568124109, 
    -0.122346317369298, -0.171442452160079, 0.186031807597346, 
    0.455553000877974, 0.321725196219469, 0.0577715045311525, 
    -0.13794021023411, -0.159282389017574, 0.535410047671913, 
    0.132800237852512, -0.109450111264203, 0.27963115647215, 
    0.449799820694707, -0.161772309321115, 0.762707210750822, 
    0.583387957989321, -0.0442446513099796, -0.0903463159744664, 
    0.815533416476633, 0.849132079510247, 0.563667072307179, 
    0.301889278214461, 0.111449591392726, 0.03353294256394, 
    0.372076674070974, 0.24218869075134, 0.0139665728465706, 
    -0.0966426769609359, 0.0742061578866359, 0.121835705247807, 
    0.000633862440864982, -0.150343433410827, 0.0329208296987834, 
    0.254504336443698, 0.0289356567821899, 0.0132864175571061, 
    0.0637342480752698, -0.0514164964367315, 0.0710308816314555, 
    0.206710258806075, 0.090186781667332, 0.00439060596566566, 
    0.0458850182382142, -0.0875611570502464, -0.017952708903918, 
    -0.204843914109746, -0.0841680425308467, 0.00372635604713546, 
    -0.0352202025091419, 0.116515928626579, -0.12461492690225, 
    0.0442348968089378, 0.0941782665308953, 0.0847730945000895, 
    0.154334904935138, 0.184005303709366, 0.133758354277327, 
    0.102720716625724, 0.128642678487883, 0.152701977374759, 
    0.148167352742663, 0.177605396525065, 0.165365505156041, 
    0.16037556758935, 0.177301437518839, 0.178331864932133, 
    0.157788691956892, 0.110369588766982, 0.139766936289156, 
    0.443381758002768, 0.274031529134885, -0.355489449285264, 
    0.207291645153332, 0.705278236340055, 0.236184599327357, 
    0.053003186481656, 0.178298960010036, 0.356215115691359, 
    -0.344548279266909, 0.609890527651082, 0.69920498930624, 
    0.13460029154083, 0.149157552132273, 0.135163421371335, 
    -0.0573381114507217, -0.0619582057500497, -0.0327885038075987, 
    -0.0847205806971288, -0.157414383041038, -0.0345322121022977, 
    -0.100274480371264, 0.0482572004582481, -0.104271333711976, 
    0.0800014248356987, -0.107196492041878, -0.00298321319122918, 
    -0.0303095193367642, 0.0564909390561041, -0.0265953058133607, 
    0.123292633244012, -0.0721759177257821, 0.138119366350219, 
    0.0526851192770345, -0.0307146451842761, 0.15822473863344, 
    0.214551236010064, 0.113883876516227, 0.0721480810470423, 
    -0.00984694310774348, 0.303714060964905, 0.0494504878812587, 
    -0.0500535826356541, 0.16496009202594, 0.630844558956445, 
    -0.0326957662084633, 0.0682766293070677, -0.454728972681339, 
    0.65586610038943, 0.484595810842461, 0.147844811854735, 
    -0.0332381899509231, 0.367795268523944, 0.302787771040044, 
    0.117501551310271, 0.0764483669754623, -0.0524504227139548, 
    0.146199599133384, 0.0316610647197627, 0.591653475413645, 
    0.16479529153629, -0.114496206846941,
  0.0122752455786455, 0.0643819737521317, 0.0626698346779502, 
    0.0449095775182297, 0.0501428876023591, 0.106631337914983, 
    0.0997862630932436, 0.0248766438579882, 0.128114819250186, 
    0.131093230248716, 0.116661628546886, 0.195795248596553, 
    -0.19285435122812, 0.72154538074135, 0.143852731556459, 
    -0.101775951605138, -0.198482874461995, 0.629434066996046, 
    0.423929909833196, 0.162111869560533, -0.284589694593464, 
    0.242891072479928, 0.403219755619484, 0.00606554847012135, 
    -0.012222357200898, -0.0737965119359641, -0.067216633995072, 
    0.0152041895512482, 0.643398226336237, 0.054651222825567, 
    -0.299914074882586, -0.134090458716914, -0.288215764283363, 
    -0.0230995565509641, -0.332485758977642, -0.0831128202034203, 
    -0.295439035315302, -0.212008909683566, -0.0436629731921387, 
    -0.267782530028646, 0.0117374890785953, 0.0982618410614475, 
    0.114125389424366, 0.119861429417523, 0.126967812277817, 
    0.120807514035484, 0.124289957892123, 0.125038854144876, 
    0.107880471907107, 0.0949439286539985, 0.115418520694018, 
    0.117049625674248, 0.122927119705938, 0.141307104360911, 
    0.154684097124942, 0.113851492796435, 0.0846125046351497, 
    0.162235113430101, 0.157478420066882, 0.154907194056849, 
    0.174628327076996, -0.134611306539157, 0.146990880087677, 
    0.467966383233927, 0.159592447289656, -0.0553303393402289, 
    -0.0132735557786318, 0.46827576167371, 0.249305618466943, 
    0.0826187649261046, 0.18368707417077, -0.0330458583555662, 
    0.410944967198812, 0.586903844649272, 0.0104454193578192, 
    0.023450608659891, 0.42529943512586, -0.330917209797016, 
    0.295879555087881, 0.263580626141146, 0.00331749288169965, 
    0.0714412625172482, -0.0480731894588632, 0.0671637330276988, 
    -0.0181188498937384, 0.0941352329914471, -0.359412185194655, 
    0.0519226407527179, -0.261846993973363, -0.171030019797592, 
    -0.00794789375828409, 0.0478681601911929, 0.140079133215844, 
    0.184784113329889, 0.209041271208635, 0.171623749567048, 
    0.13003831169861, 0.171788807119997, 0.218485250886926, 
    0.203038488026013, 0.198730950894044, 0.172683922282843, 
    0.163421410287922, 0.228608560458998, 0.27860994996368, 
    0.211759443312286, 0.13928894850077, 0.239464854914261, 
    0.346004741764029, 0.220252834772761, 0.0789161351277567, 
    0.133761248152983, 0.392582566026705, 0.267698548337536, 
    0.116915553260342, 0.158469353355723, 0.286417167418616, 
    0.43846239911136, 0.293684488572074, 0.0263320498545014, 
    0.590008696949211, 0.416496098110679, -0.167050626913737, 
    0.195499334894443, 0.838742780706124, -0.0785602556889251, 
    -0.114188425200255, 0.0836432755321693, 0.593389970765494, 
    -0.0479908941427112, -0.071771584783638, -0.179622631272436, 
    0.0461607744099622, -0.108141779692777, 0.0302096003015499, 
    -0.137434200797297, 0.0447986779638049, -0.176361512745383, 
    0.0307834365457794, -0.21340346455835, -0.0101715071821228, 
    0.0536972436852234, 0.0890004566166217, 0.172895018772766, 
    0.202828572001853, 0.123447010631151, 0.0846659916414924, 
    0.167873110222477, 0.165317320724342, 0.103238155152605, 
    0.149789345454193, 0.156045891295123, 0.132558502898305, 
    0.243732090572767, 0.306255475396704, 0.175719770232853, 
    0.0775131600261725, 0.24381788521736, 0.247216071369624, 
    0.240733195351237, 0.495436658903601, 0.196352373524117, 
    -0.0978098475948179, -0.162116904873503, 0.505028656620984, 
    0.388387939728376, 0.273202601158625, 0.0829575028400729, 
    -0.200428421074376, -0.16581004491537, 0.57839918588102, 
    0.165777667838739, 0.177077052235756, -0.0149967401724387, 
    0.519231652871114, 0.039232267810544, -0.280762082128651, 
    0.184403383190113, 0.517434002395331, -0.15173641474917, 
    -0.0900487373669692, -0.150955551138929, -0.0913123946947002, 
    -0.00354993793352666, -0.0827209639964048, -0.000261570483541862, 
    -0.120337228760135, -0.131807419745598, -0.0297983198595137, 
    -0.0860906928826335, -0.0580241330394619, 0.0232069463462665, 
    -0.151762576376756, -0.0423572084089866, -0.00168370645323854, 
    -0.107883050561088, -0.00361799598254359, 0.04522452758167, 
    0.102106579195604, -0.149789329310786, 0.0694010248960597, 
    0.231734246163265, 0.0384398399341253, 0.0263491215357979, 
    0.230228584376473, 0.435674360181396, 0.188201766850771, 
    -0.212052823873152, 0.142111465505481, 0.555208406160348, 
    0.100585773832941, 0.01451605172753, -0.338644265505288, 
    0.305129082400048, 0.501777799377055, 0.435670970406524, 
    0.563999373039009, 0.363656546596344, 0.130539219428813, 
    0.845963707527248, 0.298939727731455, 0.0636880966510761, 
    0.0133115148856485, -0.0676598675347068, -0.101989748782822, 
    -0.0267533873602211, 0.0808553049292991, 0.20190946445542, 
    0.135511421985898, 0.0285077194920497, 0.00365690499514289, 
    0.0721975340333795, -0.0781370788665898, -0.0672212938195656, 
    -0.0556182585879886, -0.106168981670178, -0.0621756995282412, 
    -0.0342743155353866, -0.0417051331177236, -0.0582610815241697, 
    -0.0941170295043055, -0.0564347187602774, -0.119328573219953, 
    -0.0689359282142765, -0.028938695907718, -0.127791587383651, 
    0.00465259811733182, -0.0151360888718333, 0.0222829698391031, 
    -0.0987654214798638, 0.00941402693570452, 0.0653815475792499, 
    0.088220034301874, 0.126763823166386, 0.149609264134118, 
    0.118961926374983, 0.10741315180359, 0.124511924431529, 
    0.055220916682381, 0.145158294590639, 0.409263719356455, 
    0.123275359913407, -0.0323193592324687, -0.202398410693518, 
    0.231932276109457, 0.570032749723535, 0.245585641746209, 
    -0.0859239265775565, 0.303055463973177, 0.386458884104549, 
    0.218272434129838, 0.215531002750247, 0.0899336118450987, 
    0.256374727500873, 0.697896622562215, 0.292622785185174, 
    0.122774045759025, -0.192537263700337, 0.363494998149295, 
    0.0721810787727793, -0.348693665823852, 0.112667152794158, 
    -0.40778504745134, -0.161747553698525, -0.10855365623067, 
    -0.251795989770673, 0.0608037195954451, -0.217957413241163, 
    0.0920168248843866, -0.275299500719498, 0.0316641061638321, 
    0.0175115939869396, 0.0600835166138746, -0.0721840557214328, 
    0.0440727416760584, 0.000772793091989341, 0.0547209354875987, 
    0.0466162907569719, 0.0695919239535237, -0.0961094975121307, 
    0.0324891893689316, 0.0291181862405604, 0.0683579433371559, 
    0.0967961180022657, 0.086242578458552, 0.0651983569348269, 
    0.062506249066585, 0.136953438500409, 0.0995747900560276, 
    -0.072529259314629, 0.139030217096531, 0.327809522855086, 
    0.140498809995846, -0.0965094579905651, 0.368834823898884, 
    0.394420207649927, 0.132869441417748, 0.0288526224095884, 
    -0.0389152133863172, -0.155950592934156, 0.401324742266902, 
    0.6419843579503, 0.0744385766376966, -0.158864961089049, 
    -0.0471316308882186, 0.57744848992616, 0.109461228877689, 
    0.132601655175488, -0.22131950395892, 0.406281178594293, 
    0.266096557557561, 0.0278940240483287, -0.142546222250568, 
    0.0647969898036122, 0.0918083906770302, 0.100467082725168, 
    0.003091973476451, -0.230733965750197, -0.0871448258261464, 
    -0.196214635696761, 0.110282404843717, -0.211145458137075, 
    0.150527279786266, -0.0923047941618606, 0.184586800491235, 
    -0.0807789213975804, 0.16438580596111, -0.149984804370073, 
    0.12927840541774, -0.152802011416014, 0.138201370797473, 
    0.00451283843534457, 0.0346152456176672, 0.0374011230467145, 
    0.0550563436504957, 0.0151968749327087, 0.0467151583640493, 
    0.0246622196737138, 0.0285011935893393, -0.0432350848092018,
  0.0680190379040766, 0.422009108995438, 1.12596474601914, 0.119775180374594, 
    0.133128523570986, -0.545727887340593, -0.0840277245973069, 
    0.851390575043644, 0.334871602013777, 0.0526423096849831, 
    0.147753826401092, 0.267793198191155, 0.0240110413901014, 
    -0.0354647878176723, -0.0547272208524256, 0.188294906520363, 
    0.199932119006449, 0.0752085058045229, -0.0674462247159919, 
    0.0843168502120632, 0.197906902939268, 0.093159190408844, 
    0.00423752268486022, 0.165665166756422, 0.103082717523523, 
    0.022244380479186, 0.070067943759601, 0.143320102113714, 
    0.0320221972079175, -0.00251638990417341, 0.233941952521826, 
    0.169111365600276, 0.0806577109853042, 0.0507612896711296, 
    0.124302252734187, 0.102214759756754, 0.09618178871381, 
    0.211358523756757, 0.188718184223269, 0.0868895312791797, 
    0.0154013513098778, 0.0590547106299836, 0.00339715313513961, 
    0.0443620694278066, -0.00967388431116689, 0.0266412437469025, 
    -0.0432480484090541, -0.00654549015721753, 0.0293258424894298, 
    -0.0307298391688786, 0.0374939651796314, 0.125045993222648, 
    0.0564439606076098, 0.14858328579903, 0.309578261997928, 
    0.174309305396377, 0.0664830831292565, -0.072700877057852, 
    0.0979973812889566, 0.0277096175919936, 0.638527809098744, 
    0.448920957525966, -0.0138599958606774, 0.562210605917361, 
    0.467913953963164, 0.0842941057824602, 0.416423643136529, 
    0.650862445556133, 0.12234164109494, -0.110139817923392, 
    0.153878919959483, 0.241134585685891, -0.0817951368888186, 
    -0.100195024601633, -0.00593206870882622, -0.0347604306560108, 
    -0.0113263688144893, 0.0246509047125324, -0.25767408410703, 
    0.105056684902733, -0.356641423193562, 0.0386618116029689, 
    -0.292791362512775, -0.110567725085078, -0.155842463924026, 
    -0.00432620451867921, -0.271072091318991, 0.0330186937720113, 
    -0.488311867284764, -0.135801028536477, -0.0559147477372521, 
    0.0507059116179552, 0.0190359680550824, 0.0538846812319704, 
    0.0966612700931204, 0.0666892871207466, 0.0698114454975442, 
    0.057920999708683, 0.0312992093267522, 0.00916102479092398, 
    0.154045720547931, 0.0823373871818079, 0.218670699515592, 
    0.424321721652177, 0.203725296563701, 0.00844806258495186, 
    0.0531366888978077, 0.590678606021266, 0.065427527283515, 
    -0.0251901929747365, -0.176955385683248, 0.224824662921943, 
    0.540747720354611, -0.016718151937677, 0.339670163501856, 
    1.11944342208853, 0.189558526690584, -0.0325541748784037, 
    0.0914020043289007, 0.667487529032721, 0.127284083899185, 
    0.0487322154267046, 0.066694672383424, 0.105870676080397, 
    0.117531917638387, 0.0712016751131042, 0.0628355206248632, 
    0.111450903410332, 0.0940908770706819, 0.0673728789526964, 
    0.158063810974602, 0.0884396790439013, 0.0441981306887391, 
    0.264683405133666, 0.291399880382321, 0.145695715351021, 
    0.0747761979843366, 0.23636765736553, 0.327879471738447, 
    0.263673358657352, 0.253509808181314, 0.246725929498416, 
    0.170296398360158, 0.182086319499995, 0.457747977181396, 
    0.43412018197847, 0.208797105255854, 0.24202807694787, 0.538620106104805, 
    0.302414201480317, 0.0416339259024904, 0.0336585320159943, 
    0.509727594188823, 0.346559215330621, 0.15413151528546, 
    0.116796630698151, -0.159623027855757, 0.52489611430145, 
    0.346712837797071, 0.0869750123484764, 0.172634095247867, 
    0.172487726384577, 0.569417025023211, 0.390132444639077, 
    -0.04444331333229, -0.0516262166115418, 0.0036097097676364, 
    0.0923402911191191, 0.451506969984038, -0.0119791291582034, 
    -0.0779385830342401, -0.228281654404666, 0.0398315301634509, 
    0.00885402438878362, 0.160941157327599, -0.22520710243878, 
    0.230658981879817, -0.341924511132548, 0.0495233242853395, 
    -0.2520711992314, 0.004800851153168, 0.128128563355099, 
    0.0128056044959839, 0.0296354745049969, 0.0963178873095257, 
    0.129101074889017, 0.107907974081365, 0.078975097123615, 
    -0.0561403679324332, 0.032527082865554, 0.030562286050436, 
    0.0240168177450699, 0.0231934265904425, 0.0239397684673183, 
    0.041271597106655, 0.0309613794181473, 0.0273966571048099, 
    0.0479650310375279, -0.038819847786762, 0.0135310335418605, 
    0.373669708596521, 0.137031544994836, 0.168073370650801, 
    -0.188059524892276, 0.278494522455015, 0.302817984118434, 
    0.576064159172859, 0.304186146664165, -0.298454042331724, 
    0.174327327550504, 0.853980789578973, -0.0794143008645161, 
    0.242773855296039, 0.986787897355565, 0.425450169637055, 
    0.0988635444672856, -0.0614763755549964, -0.487366736192175, 
    0.332411490565251, 0.627764529957561, 0.17169343688235, 
    0.0648357796605159, 0.00047326214932443, 0.26929330728667, 
    0.0357393667807723, -0.0854473259619431, -0.0576248405049931, 
    -0.0127840932878098, -0.0407498088551661, -0.0615917406008165, 
    0.247679529990213, -0.0186224901428287, 0.0172847475293424, 
    0.0749882772576048, -0.0585220770085794, -0.00131213949921295, 
    0.0446445635738959, 0.0733516512249551, 0.0969443370346925, 
    0.0237888827668069, -0.0210981376843606, -0.00186404953640526, 
    0.00460894716043556, -0.0574572910105083, -0.0269891746615381, 
    -0.0343344500045622, -0.00859488455901584, -0.0298456811759978, 
    0.0257579012797843, -0.00271678013404628, 0.0630429755033245, 
    -0.00277140241735961, 0.0307200641159634, 0.0239042987323702, 
    0.0376361609729686, 0.0160685594199154, 0.0327356801864889, 
    0.0331459646927028, 0.0364657530901664, -0.028229361985106, 
    0.0482263667513929, 0.0814313046559493, 0.0898387467656795, 
    0.131364302439893, 0.152214128121779, 0.0786303097290873, 
    0.0885316312062858, 0.335581284798058, 0.00485884137481682, 
    -0.22195627747825, 0.0185967601345113, 0.511108514171996, 
    -0.00567299406146088, 0.0753150157820069, -0.366230526744234, 
    0.516102107856798, 0.365864500821539, 0.174107324848145, 
    0.753425016624541, 0.406592932042297, 0.056521357211761, 
    0.246197791938624, 0.383597533855447, 0.073573585462974, 
    0.595882918280965, 0.471433733833098, 0.0736913196445302, 
    0.605657666869141, 0.521017673651897, 0.0110492324421677, 
    -0.0786857952195647, -0.0241750984024676, -0.0469591057241098, 
    -0.043668467202231, -0.0209117411756565, -0.0472821393088761, 
    -0.0713977908885429, 0.0481275103025422, 0.118964894251438, 
    -0.138373133543122, 0.0620363846566213, 0.14495387677235, 
    0.315290281021528, 0.427979576391284, 0.142353603923869, 
    -0.20578515019549, 0.44087019215939, 0.545649244955985, 
    0.467587087060214, 0.214357722502638, -0.260302463944936, 
    0.164545906531553, 0.243426850648677, 0.0660694346381816, 
    0.77467885931828, 0.640777354959182, 0.519534426175667, 
    0.659652573668935, 0.107017671117703, -0.381467426861851, 
    0.0548608288002422, -0.220829502556008, 0.164153593982847, 
    -0.332253645440348, -0.02049839730032, -0.206696441044317, 
    -0.182474836319952, 0.0168485565250114, -0.313606145578018, 
    -0.0594380688572525, -0.0108483629979977, 0.127694671819329, 
    0.14438965730637, 0.146956390266988, 0.0637968181822699, 
    0.132880373727316, 0.0528805458951293, 0.111810980559907, 
    0.0090723040951616, 0.0735863603680703, 0.0235772354774449, 
    0.0652141612287331, 0.00403564220046218, 0.0597685895600244, 
    -0.0144940649859147, 0.036067114905682, -0.0180580026181483, 
    0.0247987901714841, 0.0838468120215569, -0.106760288326605, 
    0.184314403131297, 0.228918494777911, 0.00233275515249951, 
    0.292291327976752, 0.30475440719687, 0.00176777444817142, 
    0.081437581538182, 0.512813499024975, 0.207929322815973, 
    0.0916131693336684,
  -0.348227370656473, -0.0293135396871212, -0.192077036412806, 
    -0.15579531940025, -0.140553891506271, -0.165283902531802, 
    -0.0345117537292031, -0.182685428290857, 0.0838569593689557, 
    -0.204515096246962, 0.109343436616032, 0.0857271237591017, 
    0.0489398340351629, 0.250264459702554, 0.289876968571587, 
    0.143156121836957, 0.0791055887440629, 0.328491360976376, 
    0.290095314362266, 0.108837938790274, 0.0469573261809865, 
    -0.12993272535737, 0.281120246115736, 0.488915622996364, 
    0.284761513188228, 0.142001884709619, 0.0690300182655812, 
    -0.0832594336706185, 0.07532373167834, 0.478380156556333, 
    0.4125791716361, 0.264503380737282, 0.18953269092814, 0.166173181061806, 
    0.148436601469599, 0.224514165976889, 0.429195183194906, 
    0.345667501935324, 0.125907421851099, 0.103235487996682, 
    0.503464816522339, 0.270746938735713, 0.0131555988495516, 
    0.158246404762152, 0.460599117848803, 0.153687505172024, 
    -0.121261569412018, 0.285267625162524, 0.455198138096527, 
    0.100221992136064, -0.121263943290402, -0.0147956165820244, 
    0.570894258864802, 0.253398325147242, -0.0513853432146022, 
    0.340298621270978, 0.382880527540866, 0.0915336439783469, 
    0.339774805144451, 0.498434418888014, -0.00204524880572118, 
    -0.0260614717860014, -0.0317809806325688, -0.0514399401549873, 
    -0.0620090587412544, 0.0538425837649448, -0.0926369168326179, 
    0.0507616520160582, -0.0333078195970452, -0.0689799735995864, 
    0.0389865380383979, -0.167534841091193, 0.054504117204589, 
    -0.081876793505316, 0.0292861099422208, -0.137913357169992, 
    0.0253878481037554, -0.150907174294005, -0.0172113465299812, 
    -0.188602675723644, -0.0555396387704101, 0.0148209400137479, 
    0.150238256377131, 0.0848514592203573, -0.024067059617011, 
    0.0431314822166277, 0.260767035499749, 0.102162488331099, 
    0.0114915834425136, -0.0575396671054911, 0.146718463159658, 
    0.0842491336804194, 0.778997246775862, 0.549690811421839, 
    0.524606562584935, 0.426021418505948, -0.157019437299217, 
    0.14215550636957, 0.681717077138439, 0.209583584633624, 
    -0.13017157806292, 0.0442145717820532, 0.45113644190352, 
    0.213663622406122, 0.11269600833242, 0.197033682628848, 
    -0.095506900828071, 0.181630710313628, 0.644124524214822, 
    -0.025148211095888, -0.125935721935671, -0.237049750672324, 
    -0.0483027280798444, 0.148610219491603, -0.105178575159372, 
    -0.146611167673714, -0.0298431480937371, 0.0359501866842918, 
    0.0474832451315915, 0.0289216809259117, -0.0331446499692567, 
    0.0133833812352499, -0.251627595212482, -0.0269119720325048, 
    -0.0742955859863809, -0.14734575085091, 0.0460583725979558, 
    -0.0435771467930824, 0.0865547087157762, -0.138218151865678, 
    0.0345637873389581, 0.0693689596713282, 0.0675928075662393, 
    0.108721188038391, 0.122471624230805, 0.0856641731884486, 
    0.0752581456705181, 0.123015936875349, 0.124018298298427, 
    0.0585557732382329, 0.0288821929977611, 0.0876066966466324, 
    0.337620330239933, 0.234480443952511, 0.0905618500846224, 
    0.137357188465248, 0.245834225480601, 0.496823855227845, 
    0.278117229695202, -0.366918922861326, 0.287850981804693, 
    0.714617348791484, 0.0465007230360907, -0.0985036592932094, 
    -0.240166251492272, 0.198515749984714, 0.938941724962745, 
    -0.0709723898502431, -0.179829623238142, 0.098787528228787, 
    -0.330076786811443, -0.150734998605467, -0.227858386306509, 
    -0.221790379280699, -0.13338567896427, -0.248335281331487, 
    -0.115302048602269, -0.189048909197634, -0.159891516558671, 
    -0.121696951205037, -0.0123409791232317, 0.0648459628604477, 
    0.0237870459114382, 0.0151494544451744, -0.0803925012817904, 
    0.0118384746875543, 0.0150909157084172, 0.0237064361401763, 
    0.200632925202411, -0.0791330977558337, 0.017481750589854, 
    0.060302425797598, 0.0718224308576905, 0.0902276971682917, 
    0.106175139091535, 0.0831332472317374, 0.0753300946264417, 
    0.107404971082212, 0.0926008457186846, 0.0444888510657442, 
    0.121047261393476, 0.159742445159611, 0.137898901436014, 
    0.16074052311827, 0.236736149592212, 0.237295579436266, 
    0.224021916909746, 0.189693834445887, 0.0807902925241688, 
    0.0347880758767156, 0.373838965035646, 0.439788470338784, 
    0.260208187548339, 0.148999850119519, 0.344405454109337, 
    0.272345724642359, -0.205756862410132, 0.360527464722412, 
    0.763995203015014, 0.490756593511231, 0.0892635430713749, 
    -0.223876594936388, 0.048560871046161, -0.135580483326039, 
    0.528689493126478, 0.392002273655902, -0.00670512530309748, 
    0.228483892872217, 0.654980255793255, -0.00607074951801465, 
    -0.0152550502259844, -0.130743821125469, 0.261102002999862, 
    -0.321432515945236, 0.168732756207908, -0.228498761680385, 
    0.172396447184458, -0.200919557382481, 0.188496059677208, 
    -0.222599053414918, 0.114786493223771, 0.0499654825448281, 
    0.113250153587417, 0.0149240170022546, 0.0696842003067845, 
    0.0988457428094724, 0.0881304649042491, -0.0521858469363193, 
    0.0654709692769907, -0.0300120868042001, -0.06950976137811, 
    -0.028816352283913, -0.00126694912407825, -0.00610320461140133, 
    0.103939856692372, -0.0277553960961828, 0.0404857219801507, 
    -0.0436873448895164, 0.0253095045920901, -0.0879992839300955, 
    -0.00217403671183919, 0.0433613336969452, 0.0616258966371937, 
    0.0560153095809938, 0.0478545324608806, 0.0571506896862517, 
    0.0855845174455298, 0.0716848026284994, -0.0253313346748454, 
    0.0286653536244259, 0.360961009970835, 0.134422151381289, 
    -0.0541685000918901, 0.42618340467962, 0.279083044298902, 
    0.131530545305465, 0.354176585995039, 0.286952213088868, 
    0.359179571423673, 0.401849694660867, 0.135349954779424, 
    -0.387972418552738, 0.326063262467698, 0.66852312075366, 
    0.332394995311752, 0.113571899147291, -0.294546959099995, 
    -0.211767249209769, 0.530186413191577, 0.503135640990231, 
    0.0875982344625568, -0.0205078819725799, -0.141567528034877, 
    0.409747184843546, 0.184337288946128, 0.0836345719357531, 
    0.0922514290624783, -0.00986142207786318, 0.168722053829431, 
    -0.171126608263296, -0.413730757178241, 0.0643959155736953, 
    -0.275673053812684, -0.136469189872347, -0.160609458045279, 
    -0.162866136276708, -0.105752396238244, -0.172066122856219, 
    -0.0406230820930913, -0.192304978526925, 0.0373704248806812, 
    0.0650560762981454, 0.0597451484778932, 0.119419536264167, 
    0.106538842600705, 0.0553405453167992, 0.072672070695088, 
    0.236801658158662, 0.232657751556585, -0.123890365212772, 
    0.525624039326634, 0.229183218194936, 0.0581230283555498, 
    -0.265876542521961, 0.189258012417742, 0.592866523997742, 
    0.190056704531481, 0.0363192744579435, 0.13985528380375, 
    -0.12817445308285, 0.164428259508455, 0.610715146050765, 
    0.350517501962147, 0.142573857834286, -0.182256150391017, 
    0.261462692012002, 0.274903768770379, 0.0215685990267173, 
    0.410114877906104, 0.435730957759753, 0.11453582490193, 
    0.0606063149162714, 0.0635798757039816, 0.068814996871536, 
    0.0781803984061837, 0.0559282962390946, 0.0195406618700809, 
    0.163354272800964, 0.0870727466770442, 0.0351330504545482, 
    -0.141638106823006, 0.539402055741718, 0.105067484711909, 
    -0.0985325330898957, 0.032913128798246, 0.425203864537745, 
    0.155810423978822, 0.299405987872737, 0.472498623641544, 
    -0.284910067273139, 0.611383909033614, 0.811378431746445, 
    0.0258959989240944, 0.158677353437559, -0.48370793006217, 
    -0.263351826421494, 0.599820986098094, 0.637678043053525, 
    -0.0357716873418389, -0.219258488429245,
  0.161219735893339, 0.073623546845518, -0.127276339098808, 
    -0.203873835729673, 0.283721669706864, 0.806158322687324, 
    0.126098626363259, -0.304213253061025, 0.0784475237706284, 
    0.636996341089864, 0.0988909222781593, 0.115771916515869, 
    -0.352469570222051, 0.172918025543008, 0.586032021550488, 
    0.384504414163912, 0.144166632957278, 0.023599959794654, 
    -0.2607168825949, 0.107458100145692, 0.392867917951226, 
    0.387496196623817, 0.24588298715733, 0.127577515070263, 
    0.0721260751467733, 0.0462126860573989, 0.0460984682123707, 
    0.0612353012623284, 0.117902632621703, 0.152867919768415, 
    -0.108803195818178, 0.119301314370862, 0.472770578593326, 
    0.251196660509693, 0.0618789843124331, 0.536346620045033, 
    0.256663125870751, 0.0184311798477837, 0.268576778409018, 
    0.397840528862627, 0.166978227701684, 0.100243954742728, 
    0.00657994232887523, -0.219844325820898, 0.792752373064016, 
    0.221488421314155, -0.167007326306011, 0.378728325423558, 
    0.460491901761335, 0.0259446047965514, -0.0797736391636454, 
    -0.0284312820707801, -0.0467326319134561, -0.054971932249451, 
    -0.00284032150757577, -0.0626816905302787, -0.0144009174363395, 
    -0.0414563343112987, 0.0195022565618458, -0.125378657908748, 
    0.0714298470892178, 0.277529846240873, 0.112079669354201, 
    -0.149987214327913, 0.303117942717463, 0.354587504349842, 
    0.0888368934875493, 0.00452248475280337, -0.168626385438359, 
    -0.084034782588901, 0.622534274957032, 0.0179956222075809, 
    -0.142211322088592, 0.16802593805122, -0.174666645506593, 
    0.202838894485101, 0.872972538790011, 0.238570114929678, 
    0.107075121270097, 0.168583307359143, -0.0659863719143852, 
    -0.220065265850002, 0.124104681807542, -0.116016110878596, 
    0.0699206302454395, -0.142146681109275, 0.00653557590832669, 
    -0.0384302612719443, 0.0657714535687445, -0.25677506093672, 
    0.0331859506469752, 0.0987516521737358, 0.117836078127796, 
    0.186816339256727, 0.191495727417745, 0.115909957724621, 
    0.0929075890997269, 0.240398942604612, 0.180907223560803, 
    0.0269393325434771, 0.0555124034853384, 0.107248097622275, 
    0.265682035492297, 0.488014496886433, 0.26498433563805, 
    0.316719727176748, 0.740533693069584, 0.138670883141806, 
    -0.0359263606908301, -0.0093721167283187, -0.288491869568233, 
    0.707103759636762, 0.467645598049875, 0.0495763068812195, 
    -0.636738211828148, 0.562614570005331, 1.18412110494279, 
    0.214216326257578, -0.139077442310442, 0.304862440126081, 
    0.392858432034822, -0.00423153056615129, -0.353373571835672, 
    0.414483943719081, 0.433783590387412, 0.0586055053722217, 
    -0.224128369103834, 0.151751923209299, 0.249311022040751, 
    0.00726581386967854, -0.123459894858718, -0.10634557750048, 
    -0.167455917513476, -0.0878943012602577, -0.108453612676315, 
    -0.0857479221775581, 0.0267336707916312, -0.0785385087057539, 
    -0.0244187063430066, -0.196322262385194, -0.0289342708550547, 
    0.0275248572372332, 0.166428242249438, 0.222244676095909, 
    0.123952543887744, 0.0355067715579914, 0.154296387833991, 
    0.222703707064097, 0.15782295446989, 0.13251227734738, 0.189509983047502, 
    0.203721405202104, 0.18672911541665, 0.174576543071219, 
    0.175001409330836, 0.167177637422349, 0.127806807202562, 
    0.13522392952353, 0.290220819154483, 0.172956426047586, 
    -0.066658148598231, 0.0224509296384156, 0.444364201765908, 
    0.387912541512404, 0.0979538423101957, -0.18020422267644, 
    -0.20757637532617, 0.329997950619029, 0.490686967848295, 
    0.278564857866572, 0.308889449144667, 0.527590325001131, 
    -0.00574529345187451, -0.147622742846535, 0.0991586596309518, 
    0.355878637979916, 0.0112047843417687, 0.577715582717734, 
    0.465932031998133, 0.0317205428252951, -0.0909763933316576, 
    0.0687600897459102, -0.165057028789684, 0.00556533416116919, 
    -0.21817403896716, -0.106015543036072, -0.0289168461333806, 
    -0.13590206914205, 0.0512958583965364, -0.159732284598651, 
    0.0459276503970292, 0.0344441947797433, 0.0889573310238486, 
    0.195562359302494, 0.230993887019593, 0.246651650110969, 
    0.172658719639667, -0.103115945997724, 0.407553528618452, 
    0.2612727147492, 0.137446674029907, 0.218510218745114, 0.169927580704992, 
    0.0666236671286467, 1.22571330263766, 0.283491700659346, 
    -0.280655250005112, 0.546387599365536, 0.536587730023008, 
    -0.189899341085385, -0.0797490451467972, -0.0319196055029912, 
    0.0396735086829752, 0.040472064295411, 0.309981003338281, 
    -0.12804728479495, -0.0956249555836975, 0.0663118521810395, 
    -0.0217030396245766, -0.179216306425268, -0.186452752208668, 
    -0.068012973005516, -0.130262193729143, -0.166317670592746, 
    0.079158176557897, -0.171655265233163, -0.0339165230082397, 
    0.0109457011937969, 0.0779844452639981, -0.207570131282956, 
    -0.0340161650766157, 0.256960227844055, 0.154471630127581, 
    0.0585605644911275, 0.043819673463618, -0.264547657740625, 
    0.274616425080432, 0.513431388316365, -0.180928478049705, 
    -0.117112353315155, -0.196459409409997, 0.644183895227082, 
    0.126215253039684, -0.183866671724783, 0.456544839213137, 
    0.401465365779309, -0.277541217189555, -0.214979058360218, 
    0.00628639599854321, 0.595015709746059, 0.185511745781991, 
    0.245179192471925, -0.171518336907779, 0.181674062410026, 
    0.2857822287018, 0.188735123806225, 0.185817105025572, 0.16565764697519, 
    -0.0854492222730889, 0.519918406954543, 0.223652799499765, 
    0.0449163096557976, -0.186744713179671, 0.164237675420538, 
    0.374682809048084, 0.224579833204081, 0.0580734591778814, 
    -0.167274342417617, -0.0426734818283976, 0.293915355170801, 
    0.179925666213974, 0.100625509309127, 0.0851106156890137, 
    0.311668422219663, -0.014696245221872, -0.018908119545308, 
    -0.0491269522108959, -0.0112608508223952, 0.308515807632749, 
    0.096941115508075, -0.0662477231222785, 0.0383690772643449, 
    -0.0796700529155654, 0.0451117245911945, -0.0294220978576916, 
    0.0649167539714084, -0.199610536257111, 0.0107909736968077, 
    -0.235144088303619, -0.147218115797838, -0.00539555870251908, 
    0.0802149549772842, 0.0737421342593216, 0.0651895439865904, 
    0.0646037324162791, 0.0977790594232132, 0.1215123769354, 
    0.0884369525500242, 0.039253124341999, 0.027672251670483, 
    0.0956860846266821, 0.127940997705929, 0.153353264081695, 
    0.169403825303112, 0.146016373889973, 0.16555225012928, 
    0.271599122116036, 0.188138501592859, 0.0421054817626535, 
    -0.0541877869663238, 0.303000410858079, 0.312810363804998, 
    0.378884916166517, 0.404734232380906, 0.127418756425097, 
    -0.248628417550698, 0.239970694431399, 0.425470326978208, 
    0.280685213968528, 0.735121862386645, 0.412564193623782, 
    -0.0546943403568014, -0.0474143117008, 0.221734207238611, 
    0.132510387623666, -0.468907613873273, 0.0555844803053684, 
    0.516304469005381, 0.202854781227932, -0.0630227749850865, 
    -0.17259789011445, -0.331921171303658, 0.0631922946899358, 
    -0.0251570863196738, 0.108952368120725, -0.263677381277682, 
    0.0537277269558859, -0.102156049271957, 0.051286185970079, 
    -0.404645099746202, -0.0459110997505745, 0.0814489642203696, 
    0.130321936629521, 0.119293970381686, 0.154421176487909, 
    0.0948841491229494, 0.115324038339384, 0.143551330168438, 
    0.110905781704202, 0.0192325819811081, 0.0318970995736218, 
    -0.013991431409818, 0.0109304525643915, -0.00840064965722069, 
    0.00997710156311929, 0.0120105273712623, -0.00648642639431157, 
    -0.0108144593014634, -0.00150449219094392, 0.102374667965303,
  -0.0281505927047157, -0.0634737429952227, -0.00848898539635606, 
    0.173966039728438, 0.247626874804253, 0.0854375745035865, 
    -0.0351571951430287, 0.15561802836277, 0.0500225664575085, 
    -0.100865223297044, 0.0367227940853837, -0.204687571400594, 
    0.148252240179677, -0.157698031713803, 0.115288961509936, 
    -0.212140341380051, 0.104307975149372, -0.190500489959621, 
    0.0593645594570771, -0.235719530970741, 0.0257468883760686, 
    0.00286318981094615, 0.0592632256648042, 0.2399833332378, 
    0.15860649090822, 0.0190322556693976, -0.0277818639392929, 
    0.346547208599263, 0.26463137467949, 0.196386803031282, 
    -0.235281281962376, 0.45412506993586, 0.436889726028602, 
    -0.079935470529145, 0.51599282179911, 0.645067096876624, 
    0.527423652404611, 0.363369985806613, -0.214981304094732, 
    0.342846602973884, 0.420482593671492, 0.384391210687604, 0.1865619652688, 
    -0.290619640252097, 0.104253043694351, 0.437291138681358, 
    0.0881340107103531, -0.0512753308379853, 0.267983525929765, 
    0.314830170330492, -0.315791790060352, -0.235084853283334, 
    0.051266871487983, -0.0301556338024352, -0.074964862340828, 
    -0.0401326471375827, -0.116830806894837, -0.0239884054087268, 
    -0.0342245485819845, -0.161515405086623, 0.0671611533087365, 
    -0.0606726498942865, 0.133474906874442, -0.0538642091751746, 
    0.132432212669344, -0.133182564658231, 0.073658786046968, 
    -0.0604702025133013, 0.0911711719828481, -0.147908331602723, 
    0.0316698107586925, 0.0358168459742269, 0.0457822225302015, 
    0.040273604164311, 0.0477621074500126, 0.0343856942749213, 
    0.0117887111006135, 0.12532073956303, 0.0618566217501187, 
    -0.0477865717773309, -0.111290297934856, 0.196955572504504, 
    0.355557451755678, 0.20081750792107, 0.107778071566431, 
    -0.255108749370884, 0.375188026331208, 0.371008951981052, 
    -0.090881291121981, -0.135245485200524, -0.109782487248697, 
    0.163112142815501, 0.0366748587038038, 0.888137708278294, 
    0.41631529639961, 0.0289415676468118, -0.492554779852159, 
    0.567563715527498, 0.667954465791621, 0.0473188168554085, 
    -0.147630649644294, -0.180059766909871, 0.133326083824298, 
    -0.333605687858909, -0.0280047304216215, -0.276370428252973, 
    -0.225014560162531, -0.0279643087354533, -0.262120762456348, 
    -0.191374554652572, 0.0161879891984567, 0.188675379926432, 
    0.125413647947383, 0.100336844930475, 0.176433755616673, 
    0.161630659669214, 0.138778814064691, 0.151343586127258, 
    0.261876945815371, 0.233620795620212, 0.104738291860792, 
    0.0547330715474847, 0.0774220690802441, 0.0636568261363468, 
    0.0766446718071921, 0.0602605929438483, 0.0418551484907379, 
    0.10756491643859, 0.116100338233328, 0.036364151426053, 
    0.0128549714547612, -0.0259237592870874, 0.283876970956336, 
    0.255896940727132, 0.149832517289418, 0.0961689082604061, 
    0.0938516389817442, 0.489540027128199, 0.0460905765318749, 
    0.0975959941631111, -0.40265859885922, 0.115487529751015, 
    0.467488786693883, 0.49961959951202, 0.35393168818807, 0.492225952698215, 
    0.50353414267822, -0.363135157584135, 0.3560235837665, 0.78449734427623, 
    -0.0707265512484815, -0.0480365327696513, -0.0620855943987958, 
    0.0038027234089929, -0.107342136386874, -0.0330889580022827, 
    -0.145274133019089, 0.24626387916637, 0.122265245784475, 
    -0.149453498331979, -0.18698829480667, -0.00491281124556082, 
    -0.134752320533109, -0.0154016834014106, -0.14880751883635, 
    -0.0416442932474603, -0.129024729747998, -0.0769707163055899, 
    -0.11555388777688, -0.0620172094309724, -0.0283916276618627, 
    0.0247863871357617, -0.0037412901428614, -0.00941833187587775, 
    0.0373648507933376, -0.0125916606115687, 0.0299841578009003, 
    -0.00164671901488345, 0.0295455752778173, -0.00903231811921273, 
    0.0507600457307795, 0.0969430929438471, 0.093312930156221, 
    0.0956206472875092, 0.121321707477375, 0.116395947466874, 
    0.102700086551891, 0.112529375905188, 0.0900541071238022, 
    0.113996050854325, 0.194936537668922, 0.0635291547789713, 
    0.00302860773429976, 0.439600671637026, 0.253316310389907, 
    0.0654566108040653, -0.0261024467330969, 0.311702190501243, 
    0.234613678704939, 0.130412337077554, 0.460523105105077, 
    0.35601585699589, 0.18754007303559, 0.184372331962745, 
    0.0478069571285587, -0.343869453342987, 0.571770728681162, 
    0.428931404360622, 0.344716766310231, 0.400134416896146, 
    -0.0834499559558458, -0.282088238793131, 0.0103816229067534, 
    -0.183092584160087, 0.0869801389527179, -0.246951593953391, 
    0.0619347193898695, -0.217441319375604, 0.0543288469083417, 
    -0.163425474872176, 0.121314775914067, -0.0106660541722671, 
    0.0657395125758288, -0.171051416159462, 0.0120837303099923, 
    -0.173143822287394, -0.0151923677509588, -0.095634592408313, 
    0.0584630874200943, -0.296233467718505, -0.00672435029614268, 
    0.00123947701408893, 0.0253473970102575, 0.00544807112010448, 
    0.0142448648982498, -0.0115161359946205, -0.0200431422703127, 
    0.0299090080821833, 0.0198020036124803, -0.0591067903349737, 
    0.0383130573698015, 0.118243948137499, 0.126078299731939, 
    0.11077204544519, 0.0871193423214163, 0.100447405072718, 
    0.236084383967586, 0.198860091215783, 0.0337681157011249, 
    0.0594386162478312, -0.273036420231448, 0.462608334292894, 
    0.303868526102769, 0.0208827931513396, 0.438925210914276, 
    0.34989554307435, -0.042339464971448, -0.269638106517589, 
    0.571908881671185, 0.558450051737974, 0.0994581677751046, 
    -0.0929822143219018, 0.0578746585110901, 0.240620263475131, 
    0.141553333950491, 0.249398136549916, 0.0897565319372279, 
    0.762973634402872, 0.536648120904478, -0.139742473526775, 
    -0.225716319510931, -0.111150874017308, -0.153131797981075, 
    -0.168170341447115, -0.157676648290063, -0.157257270118279, 
    -0.13370844051718, -0.164604313363204, -0.0372241617276156, 
    -0.205056300719081, 0.00309902247163297, 0.079248532348036, 
    0.106843588000478, 0.13420448408209, 0.150925269056847, 
    0.095792516474039, 0.066526343495269, 0.251605882027608, 
    0.134851113663533, -0.13806039799198, 0.218345035307355, 
    0.458275103823928, -0.0252490849348981, 0.327627907946475, 
    0.614177921333372, 0.301928864486667, 0.177014439705889, 
    0.0272334563512595, -0.0438199094633521, 0.340623984059426, 
    -0.0939599058636542, 0.345380944979301, 1.01479764393791, 
    0.0999340363466804, -0.0914850144774824, 0.0631831415299996, 
    0.756649363929403, 0.0148129755848037, 0.326833288692446, 
    0.959965588491361, 0.0770123600878486, 0.0111834391671689, 
    -0.00153333990112906, 0.0194591819707871, -0.00650031700215774, 
    0.00445883636322186, 0.00419222997593197, 0.0229639146491753, 
    0.0412378636405009, 0.0148740196975888, -0.0383879282210491, 
    0.0186324265899227, 0.443752796576081, 0.120506329955198, 
    0.0699024056374138, -0.201460980178896, 0.234458952626884, 
    0.450886867311874, 0.15603701965186, -0.163266624593527, 
    -0.0716024181808478, 0.469806041642182, 0.455429378096633, 
    0.071392947684986, -0.0421980814002743, -0.171778396716102, 
    0.618057739697797, 0.162379853581158, 0.113695879475329, 
    -0.0888277463133652, 0.430635190821425, 0.385878414739648, 
    0.168082633146833, -0.17488869813898, 0.0750525952754933, 
    0.4261964128846, 0.106347208146429, -0.0201144605606529, 
    -0.135421667687985, 0.248099469836758, 0.382082913024228, 
    0.128714835606076, -0.0722323943873265, 0.0164021726249907, 
    0.121325410173948, 0.471960849426287, 0.291578419811344, 
    0.0454074396012956, 0.411770861455973, 0.252101214509819,
  -0.248957171153709, 0.183884015706578, 0.703405615228919, 
    0.214292259564205, 0.788870877359991, 0.437454667443812, 
    -0.208054058310709, -0.319948074736267, 0.162842457020961, 
    0.623031881440591, -0.204952284716283, -0.0238667972046392, 
    -0.128740204724685, -0.00122732745166117, -0.145400214032041, 
    0.00233760647542071, -0.0874061940925263, -0.0763060357126533, 
    -0.150931340186101, 0.0366710813311316, -0.0953936111503941, 
    0.158164041623027, -0.0262218809730874, 0.110472341336725, 
    -0.201090835271861, 0.0110596344479664, -0.112813248887604, 
    -0.116649485122716, 0.106418390361463, -0.133012551835895, 
    0.0603244109196531, 0.011930762512725, 0.0274151469814356, 
    0.0321568195176054, 0.0326957394714583, 0.0108590283152624, 
    0.0207921631526339, 0.0268184635418984, 0.0281791075476266, 
    0.0297234292352143, 0.034011286701467, 0.164576093904925, 
    0.151677785724675, 0.0912490133915403, 0.371772639365708, 
    0.371490258149036, 0.146560953218354, -0.192572417825235, 
    0.30490794537998, 0.413647749987255, 0.229555461008113, 
    0.242777026004691, 0.421714884675971, -0.328325395052506, 
    0.163638631903852, 0.844708171791153, 0.439736414612795, 
    0.22817296048932, 0.325246979743812, 0.560127445585416, 
    -0.225101788631247, -0.133617381308995, -0.191385125356973, 
    -0.139003165164531, -0.115975155126326, -0.154353818980121, 
    -0.00889042535774685, -0.15153219952026, 0.103089736542862, 
    -0.202043662236692, 0.0575764543937007, 0.0890755474666581, 
    0.12064217992738, 0.101532707945276, 0.13046182932944, 
    0.0729448394749426, 0.106579277656903, 0.0748256998933764, 
    0.103054959388893, 0.0760614316063408, 0.0863408070126858, 
    0.0749366968594536, 0.0816572113719844, 0.0857425717078598, 
    0.0876356957505745, 0.0728488162433518, 0.0833817605474563, 
    0.0896403819639946, 0.0514665669858255, 0.0339503758932173, 
    0.232950313551801, 0.141199669087112, 0.214817645118941, 
    0.221918068292649, 0.212610457830914, 0.516930750414672, 
    0.319272259679374, 0.0520362334798512, 0.620661101357793, 
    0.364739701677146, 0.0324301192478801, -0.166903168835547, 
    0.408609865923505, 0.664173187329388, 0.722006541758623, 
    0.383271217660463, -0.518457030337419, 0.705033160448304, 
    0.53460080066749, -0.544093024860259, -0.353657366571318, 
    -0.0693167955767187, -0.249669015870113, -0.14658820628661, 
    -0.21403724930184, -0.0228176399635146, -0.226038860613339, 
    0.0280673713643739, -0.23902878620579, 0.0331410881933266, 
    -0.0872573062372322, 0.0432614141755439, -0.0394273976267614, 
    -0.0375852327547571, 0.0684647164999545, -0.0662885526373083, 
    0.0376153869103688, -0.0287278838226848, 0.0105908679985753, 
    -0.0133240434904898, 0.0342795256632409, 0.060283767405048, 
    0.0377380150625686, 0.0498096205583066, 0.057900192141701, 
    0.0396339806144863, 0.033126829497342, 0.127355584292505, 
    0.0878224094691664, -0.100906797251411, 0.0452396026035633, 
    0.291564342254227, 0.0657768051166568, 0.254202429688818, 
    0.476514898379741, 0.149252027336568, -0.121159215088217, 
    0.391549256626028, 0.46779257484883, 0.243608391785281, 
    0.0378872819870333, -0.168588394616183, -0.27937735374013, 
    0.0709781757400134, 0.664443594518272, 0.250518899293078, 
    -0.0945408097155853, 0.427290142647296, 0.154072439818736, 
    -0.116988796470811, 0.082277242392973, -0.21170222153628, 
    0.165578480002011, -0.43579183488141, -0.0553576033576943, 
    -0.257113516984622, -0.254499098249494, -0.0155361549911256, 
    -0.240079402000027, -0.0558887315373993, -0.0260060212508093, 
    0.0593531870689462, 0.048625089613602, 0.121297697272395, 
    0.173778129936248, 0.0718575932539993, 0.104756252182067, 
    0.0832399573506323, 0.083588661569584, 0.0270734004010716, 
    0.0460841546843027, 0.0679865544002628, 0.100896997906934, 
    0.13755393639565, 0.151692270791865, 0.126948988349573, 
    0.122651633667788, 0.150269298102664, 0.133833812258957, 
    0.106739791832186, 0.132781536564684, 0.164854001121884, 
    0.163898510962015, 0.162474624291585, 0.181207186831946, 
    0.175903453481686, 0.160429115396279, 0.184212127799013, 
    0.203968860290643, 0.200576928594895, 0.16469339335001, 
    0.0185151538422633, 0.17798896743726, 0.441964528337838, 
    0.239038457153292, 0.0746077461601061, 0.129589670464635, 
    0.16055404538428, 0.229738174669199, 0.545489528079508, 
    0.367310472925117, 0.125003215219066, 0.244712924380159, 
    0.318580379760187, 0.10237146227209, -0.130265731336881, 
    0.951132169646119, 0.202609639603414, 0.0925913616051413, 
    0.012025071122771, -0.33243396472704, -0.192375030646693, 
    -0.0745618737794423, -0.277809736615742, -0.00996597873266569, 
    -0.301122899468647, -0.0666548880947163, -0.238684691602585, 
    -0.0941970912036806, -0.163085204412085, -0.010066025644859, 
    0.0727853437277554, -0.0281563736785912, 0.0106359682831795, 
    0.103822144702528, -0.0163785533846672, 0.042069905225731, 
    0.0649504002094156, 0.0637824861211049, -0.00423706419951458, 
    0.0552539083231755, 0.090871488249489, 0.0962533666653374, 
    0.138742967635307, 0.174639566861953, 0.145182823861722, 
    0.133328290466823, 0.155171279512207, 0.143135431419026, 
    0.257548577695686, 0.258165221586122, -0.00147826717652574, 
    0.0790624313023794, 0.615819805608956, 0.139687856052834, 
    -0.207563011767168, 0.21114945197581, 0.518578814839031, 
    0.0946593466827948, 0.271579118694378, -0.276918674920216, 
    0.57134569934382, 0.259330049300568, -0.00493947496919309, 
    0.00930616901167936, 0.746963105157901, 0.1931562974773, 
    -0.00389173562209325, 0.159036770534574, 0.665448830089459, 
    0.0522138218358092, 2.64035065337398e-05, -0.0501412406743379, 
    -0.0690666204037975, -0.182529034201174, 0.0952554307259447, 
    0.00410056272138597, -0.0364509521057745, 0.0580252350723748, 
    -0.0766670516547197, -0.0865914141646995, 0.0711426191224305, 
    -0.0985326846534222, 0.0717789055178161, -0.254903819482162, 
    -0.0269182604771107, -0.111485513455085, -0.0550796479180206, 
    -0.100077874810163, 0.00244270991590242, -0.0620661074223466, 
    -0.036460534408419, 0.264515073402499, 0.367760908214195, 
    -0.0149954387155527, -0.0477228239074799, -0.133398545107027, 
    -0.0659518859422892, 0.408676950089895, -0.217966460042507, 
    -0.386697495076284, -0.258640370962465, 0.312793879217508, 
    0.976747987981347, 0.335170840965907, -0.0757227598163545, 
    0.196091731099857, -0.168952398800545, 0.963164228223686, 
    -0.130647663751524, -0.197794420885212, -0.015321704659119, 
    0.0772156482080501, 0.184199391260931, 0.297662036484558, 
    0.146320434490635, 0.0283806407406273, -0.0267642701080882, 
    -0.0379991781286795, 0.197454539556112, 0.148806866149897, 
    0.0387430314673335, -0.003159450471118, -0.0390867129118074, 
    0.239458356482262, 0.123369254917643, 0.0314306674697702, 
    0.0542873020700705, 0.150918857902879, 0.0642780700595573, 
    0.0992063140812976, 0.241716140759419, 0.174388850778255, 
    0.150060540744414, 0.235905365937534, 0.135295990064602, 
    -0.0143901526219069, 0.09962311146312, 0.244717865997531, 
    0.106512022841662, 0.0158558918287325, 0.0453144722337163, 
    -0.017942919134562, 0.0148552899570419, 0.0314991753623215, 
    0.0460587625045887, -0.0401652380529021, 0.0349657954972054, 
    0.00704052224582005, -0.0495968912888473, 0.179671408452892, 
    0.0144199479630363, 0.103603689638853, 0.330311737017815, 
    0.191707329244499, 0.0976105138670401, -0.114886808086494, 
    0.290030158167526, 0.323229448216416, 0.138681944283999,
  0.0164563608162056, 0.10820145090493, 0.104790392142886, 
    0.0831309337625019, 0.139447159844965, 0.230099775901568, 
    0.243840003526823, 0.122442970083833, -0.0871300922741325, 
    0.101073413709127, 0.537498778608892, 0.100614924962805, 
    -0.152474938811673, -0.0676216111678332, 0.481391744752146, 
    0.400001099047223, 0.101538988735595, -0.166856858574087, 
    -0.104504076639472, 0.466073339927621, 0.320567053132925, 
    0.0558465035225559, -0.136022423112577, -0.0553907696430119, 
    0.106790765041689, 0.423236762530034, 0.136771072986658, 
    -0.260377288947492, -0.253900205235951, -0.150021599089357, 
    -0.0421743718277414, -0.280449135560503, 0.184846633972374, 
    -0.242077536392776, 0.169739259514176, -0.12973921854455, 
    0.13855830622336, -0.11920764376067, 0.145511528773318, 
    -0.187907665490917, 0.162430341578282, 0.0115493833643155, 
    0.0328755967943313, 0.0690056002757151, 0.103955732439276, 
    0.0527578212683585, 0.101149127492936, 0.0829246892983562, 
    0.0756536236157457, -0.0404482395366205, 0.0446678321623673, 
    0.0572623615892303, 0.0733107437407272, 0.133273078461622, 
    0.138497574014312, 0.0809122013119946, 0.0578384698809111, 
    0.231880558309349, 0.103383159875153, -0.117868293320792, 
    0.00621102306773162, 0.535979129286156, 0.134072251693131, 
    0.0389998306483662, -0.0763834519157484, 0.123992663062969, 
    0.0197351838099865, 0.872662560142389, 0.335403566187106, 
    -0.198914979923475, 0.151611854773316, 0.703618718929151, 
    0.30449552419514, 0.206912546471807, -0.235563373860887, 
    0.606664536676744, 0.566141489064145, 0.199286687454582, 
    -0.31751506752509, 0.155553800925863, 0.363249779170978, 
    0.0403347866208296, -0.00964113259036269, 0.0289279429668292, 
    -0.178489300174626, -0.224409107081094, -0.0342770378918416, 
    0.0999570985715378, -0.270683720480551, -0.108411402522828, 
    0.0177752799373396, -0.088712761407604, 0.15538541368111, 
    -0.140340127752132, 0.06487927110703, -0.15759900481263, 
    -0.0720513195207479, 0.0380509697591946, 0.0991032103123392, 
    -0.16505774574237, -0.0796085892165882, 0.00228909165047446, 
    0.534941526886414, 0.114502171123192, -0.143870734310375, 
    0.0576401384632687, 0.48232334256946, -0.0782893640164278, 
    -0.187052706944457, -0.0712048687122361, 0.57380996228606, 
    0.128590383666799, -0.324719930148096, 0.593450166266852, 
    0.53318588129245, 0.218449598782502, 0.0725952092134934, 
    -0.22029968704413, 0.0226053412292769, 0.621805033002053, 
    0.338591919237718, 0.136690043969805, 0.111401096666883, 
    0.381166856010083, 0.361488370659915, 0.155607179745131, 
    0.085694764130852, 0.305440473126223, 0.235698720803852, 
    0.0817938684435164, -0.061509450801939, 0.458388488766047, 
    0.279842782453768, 0.221334667692201, 0.259746292160268, 
    -0.212309314096661, 0.30841581081529, 0.338118058671122, 
    0.191556673293343, 0.717373506249939, 0.458510542294145, 
    0.17695159148395, 0.181962316246327, 0.146190783201199, 
    -0.0221673146041237, 0.792358366101947, 0.181896939853918, 
    -0.28284018662823, 0.32781735799933, 0.561870666963989, 
    0.155765563085948, 0.0806099507749005, 0.0713266883758753, 
    0.11023658078625, 0.119116703527733, 0.101824424340978, 
    0.163081138516147, 0.115694556327687, -0.00837963688018187, 
    -0.0292112451485413, 0.476417953256941, 0.107910214754382, 
    -0.000896047195091607, -0.114394110560068, 0.0389145342183804, 
    0.40697783296889, 0.606597053425072, 0.236816341499648, 
    -0.157628650297319, 0.18807794542026, 0.524062618861734, 
    0.145164813526627, -0.0850646921687675, -0.108048960783721, 
    0.453735011802392, 0.54223425220642, 0.0567173519483119, 
    -0.179328249093907, -0.0539582315847548, 0.488077632600277, 
    0.0578719401636683, 0.0111924220101986, -0.15878721941589, 
    0.1521284083468, 0.442738232218253, 0.143249916931182, 
    -0.0574404429497997, -0.00803436226212249, 0.439606454086494, 
    0.256280886727517, 0.126333024139609, 0.114887945390404, 
    -0.21420159525279, 0.288695893700953, 0.282087042825464, 
    0.169654775739769, 0.0837445483454147, -0.0653149388723103, 
    -0.0691377011705768, 0.38416527342532, 0.182120272468608, 
    0.06180071208342, 0.0215874720478, 0.022423166653238, 
    0.00408815291403453, -0.0284402139175052, -0.0122601783461474, 
    0.0438909584645541, -0.0376364790207136, -0.0286154075313398, 
    0.018477654721188, -0.0204860395315681, 0.0507982876366903, 
    -0.023322926770294, 0.0306385374193565, -0.0134119693078548, 
    0.0339359966485578, -0.0108456246523129, 0.0339738441589612, 
    -0.0613047805737774, 0.00534473417576945, -0.0101080024456393, 
    -0.00663187306519845, -0.00799833855731885, -0.00823067346039434, 
    -0.00586679131520949, 0.0624552281223009, 0.178832383735642, 
    -0.0880740465230735, -0.0483414657735766, 0.160699376111623, 
    0.743612311535762, 0.0609545879996153, -0.199294774922266, 
    0.0587129190772681, -0.330568022281668, 0.733860343877545, 
    0.411032448342029, 0.106828920884183, 0.261804148845565, 
    0.18336779523601, 0.19359306975675, 0.617866610062651, 0.362384848172342, 
    0.198417846753781, 0.082519079085294, -0.103685720175053, 
    -0.303067120352764, 0.569373576249583, -0.0215535552861824, 
    -0.0957473221601561, 0.0791863954262671, -0.259093371173893, 
    -0.021291714645639, -0.153114762867576, -0.128616359285904, 
    -0.0782069403368029, -0.0690745646602607, -0.21329006222683, 
    -0.0398346461409732, 0.582338276029628, -0.105530744342614, 
    0.0687209958703179, -0.431056273245594, 0.395501339437689, 
    0.680501724282727, 0.177476759652489, 0.124192803172645, 
    -0.350129311097752, 0.368033583396986, 0.409858198184932, 
    0.162344234298043, 0.0245173069177061, 0.0332279225433051, 
    0.446322381945532, 0.268272484988226, 0.0516549714770991, 
    0.375448397685261, 0.309866008758046, -0.0644119744355492, 
    -0.137567422870059, -0.120837278292348, -0.0316444959135057, 
    -0.144862157994338, -0.0260445235749763, -0.145244351363335, 
    -0.0314041102511879, -0.124184955251647, -0.0028144868829853, 
    -0.144887330737041, 0.0193652478150049, 0.05600409609046, 
    0.0712735392697596, 0.130483539629722, 0.118543753300729, 
    0.0656375214876909, 0.0801362074940963, 0.127844003546038, 
    0.168659284527533, 0.125012123593253, -0.172364888992537, 
    0.235173759940164, 0.660203274749536, 0.510036498638129, 
    0.189427713235076, -0.013414111607357, -0.0707978590239335, 
    0.822754627479963, 0.276508826005873, 0.203866300171965, 
    -0.190926203752689, 0.0709394454016258, 0.14514793667167, 
    0.522272164932378, 0.578048742083786, -0.00225260409948948, 
    -0.141234083405097, -0.271449636531372, 0.448121516065958, 
    0.340033528206725, 0.151356197684684, 0.245945027555156, 
    0.081064447757005, 0.0111036478918808, 0.00930217118011331, 
    -0.0641102944622652, 0.0461324010011809, 0.0243753319754723, 
    -0.00496578472212365, -0.0382459210767285, 0.300086848377128, 
    0.0132207814184549, 0.212757562421317, 0.448210991047059, 
    0.174788266240201, 0.0413750929141663, 0.158076391568047, 
    0.107912950605031, 0.0863562151081338, 0.480069490298989, 
    0.320701108153121, 0.140782211157572, 0.239235892459392, 
    0.282691626213446, 0.0954260035797345, 0.022432565008675, 
    -0.0137211206595884, 0.150102087252931, 0.209698385858992, 
    0.0764292574664223, -0.0399206866377233, -0.0647623816769019, 
    0.0394969678123156, -0.0625400725895866, 0.0116411900924464, 
    -0.0819802531504013, -0.00184721062184337, -0.0392053584004238, 
    0.0246669327254403, -0.0996209681837635,
  0.00429656768086629, 0.0638560973957975, 0.0992698244243614, 
    0.146157191283595, 0.148185043567382, 0.134525299776657, 
    0.16235348060735, 0.198099957421826, 0.193711005084855, 
    0.184587021385691, 0.202773787651265, 0.192693598198689, 
    0.212530975247956, 0.24031445664171, 0.215754764486378, 
    0.181625460752988, 0.202372362694751, 0.240357007480235, 
    0.219359031531207, 0.192192309430339, 0.218420379449805, 
    0.217529682258751, 0.147481203395755, 0.140141726286584, 
    0.324740902169524, 0.295307647718836, 0.119188125896816, 
    0.0465207986737775, 0.446325468393188, 0.21882486860412, 
    -0.15522219834312, 0.331387130132532, 0.529699052663293, 
    0.0325524528976844, -0.0838508328673422, -0.15214706819735, 
    0.360945888262163, 0.816768276074412, 0.176721409931553, 
    -0.154202823941475, -0.121559573601334, -0.372031522645774, 
    0.166183715691942, 0.476113784474086, 0.12158194640205, 
    -0.185073266292101, 0.0574140810613901, 0.894927634687585, 
    -0.0993782411841927, -0.104605202075395, -0.143017990047863, 
    -0.357392212327604, -0.108341848043242, -0.158522673949535, 
    -0.276599717506087, 0.0276769618103951, -0.317853364775947, 
    -0.116565612114991, -0.146107088170424, -0.26067405915957, 
    0.0183850646731213, 0.115430862130373, 0.130572002777477, 
    0.163921116408106, 0.183472421550639, 0.158003416189303, 
    0.153548125116793, 0.177702378440007, 0.180464425773836, 
    0.165698941421566, 0.168612322194444, 0.16186058008147, 
    0.155195982594358, 0.151953131939267, 0.233838602113714, 
    0.29615635941387, 0.193581551568885, 0.0905413722597077, 
    0.263044369997964, 0.342636660953244, 0.172072967104355, 
    0.111048911459237, 0.0996208019378485, 0.0941788313685452, 
    0.0974007024652678, 0.0810597163681382, 0.0849306746944057, 
    0.108001041022417, 0.0989501379362717, 0.0517267833676002, 
    0.117510619451602, 0.154975587496124, 0.109474450807145, 
    0.120724290483575, 0.228285814607175, 0.118876501800361, 
    0.33240919336773, 0.382139446997338, -0.0590151239906378, 
    -0.0755985096793537, 0.124939750194464, 0.574660640052367, 
    -0.122706588445338, 0.0191895913893732, -0.106432353566191, 
    0.652996345395032, 0.0559783652044412, -0.204160837273144, 
    0.454664569337985, 0.192018945432051, -0.256736842521176, 
    0.0656529904002691, -0.124405040065321, 0.0576119857709327, 
    0.0852009902091942, 0.00557140850773866, -0.0634309900528465, 
    0.0235196302990356, 0.14748074878608, -0.0957544731746029, 
    -0.130487883441019, -0.0145440909318465, -0.243161164030412, 
    -0.10069135694383, 0.0182906314041653, -0.152734330542879, 
    0.180928968772697, -0.0192995473452878, 0.188830726044241, 
    -0.140112430844071, 0.289732302127103, 0.242265029507611, 
    0.0618656570758507, -0.0998343695972891, -0.10784262164903, 
    0.31996023679825, 0.287456370350698, 0.180687169242926, 
    0.189498793250223, -0.313581875894116, 0.70019121166298, 
    0.415028280854355, -0.182172095731169, 0.260188905584142, 
    0.64782967569917, 0.0989772926335038, -0.221547154260079, 
    0.0185956125749869, 0.734286546679716, 0.394306529221559, 
    0.0750640868733189, 0.0975277085484287, 0.265936830407784, 
    0.282044071395043, 0.193872844639694, 0.13122057721677, 
    0.145814997171551, 0.146518689791068, 0.0487844462911061, 
    0.0755977449805173, 0.331575745531731, 0.20100337905986, 
    0.172866675415009, 0.201986755098092, -0.217967757643082, 
    0.233504544352309, 0.53147031490849, 0.0484546310599273, 
    0.0495366100629531, -0.0744684304523613, 0.263305073997623, 
    -0.0917290575443292, 0.513324581331119, 0.483424344026513, 
    0.201325873966336, 0.643073581814834, 0.461388640645831, 
    0.183951284264003, 0.219244643163566, 0.0246191319756827, 
    -0.437377119501284, 0.121797450014201, -0.317981456493822, 
    0.000278562973659066, -0.305331377466715, -0.0234982480650029, 
    -0.290437367842362, -0.196173756938571, 0.119046838218141, 
    -0.275847018863035, 0.155270591720934, 0.0379626617037486, 
    0.0497976090994634, 0.108515864689163, 0.120459784008485, 
    0.0810411665537757, 0.0938227444250891, 0.102674674747923, 
    0.107419294468196, 0.0202074706041117, 0.141169954177233, 
    0.169118724563395, 0.0508643237831349, 0.088632967587379, 
    0.321414081752393, 0.209505617289734, 0.107202913832841, 
    0.0994153721848513, 0.124477710113558, 0.114158892032599, 
    -0.177187264554564, 0.80283900019356, 0.307734562881241, 
    -0.129158208395436, 0.25539175110988, 0.577569828752532, 
    -0.00241371284180594, 0.0281834137725863, 0.956309010493614, 
    0.491732692268159, 0.0240424584271243, -0.160416527387787, 
    0.0800068238110298, 0.143672596686785, 0.138915166626461, 
    0.326016479845395, 0.177719329435173, 0.0378962842516141, 
    0.186234369299547, -0.0872708510483014, -0.356110136448159, 
    0.233479667887099, -0.322622232276326, 0.115522230398606, 
    -0.311553966466573, 0.0576638466275464, -0.351255072024557, 
    -0.0212947454434311, -0.309209764350684, -0.155042414160355, 
    -0.0370734256197938, 0.078796634050206, -0.133502840805371, 
    0.0120778790962892, -0.065282502642677, -0.0417122436085981, 
    -0.145909890844591, -0.0840938635588946, 0.016404275659277, 
    -0.183838545200799, 0.0624655503539595, 0.0624010257110025, 
    -0.0431593082702958, 0.0820683949387368, 0.168484835027439, 
    0.0382290066250272, -0.0264621965431256, 0.153279328796561, 
    0.319525180888379, -0.25302304023535, 0.134836174184816, 
    0.555863436671614, 0.41037312047126, 0.0797957362556194, 
    0.106149345710744, 0.959483094107459, 0.554644036029941, 
    0.28585335780019, 0.324176052854704, 0.379460767237713, 
    0.409366184469867, 0.100579331878512, 0.0729062007967586, 
    0.151300784376035, 0.00320977410409307, -0.153537109216586, 
    0.306953831862028, 0.176495241494796, -0.0597617149260485, 
    -0.198146809215592, -0.108980766386787, -0.287405974128328, 
    0.196204197933064, -0.17210665380709, 0.190891340439976, 
    -0.202953314695372, 0.152637129372957, -0.144335047513636, 
    0.155408778147054, -0.212370875632088, 0.0978960508013208, 
    -0.0850755097397338, 0.0134793132483388, -0.0524750473643939, 
    0.0391101507674009, -0.0994705523563, 0.0340680758596171, 
    -0.0235753518785831, 0.127979444539809, -0.0797014289135324, 
    0.226673973925375, 0.149220815582067, 0.0653337652446311, 
    0.0505103750732806, -0.171566139201304, 0.146951654748342, 
    0.301906254495447, 0.180307614911488, 0.158102491857473, 
    -0.284715148923548, 0.0767384938291603, 0.174449142127146, 
    0.711979409964481, 0.506966019829205, 0.0482858646512854, 
    0.699640260607843, 0.722696969880611, 0.186723713742864, 
    -0.0440573390262902, -0.0286338282280125, 0.607783572901413, 
    0.252268111877292, 0.0498873086940861, -0.0923665878858292, 
    0.446097116052538, 0.246543145512407, 0.0292196888677202, 
    0.0970700785780781, 0.28033313487057, 0.239931877169306, 
    0.236059430417786, 0.241441495053553, 0.235173768641682, 
    0.271555432596914, 0.0100018476920075, -0.173302544346043, 
    -0.103073892507537, 0.129377932090837, 0.185615036846655, 
    0.229272997931638, 0.14988581824253, 0.0548179222860686, 
    0.0702258466593743, 0.101589098250005, 0.00466054447008152, 
    0.068562838231221, 0.190052442890657, 0.0217711847451257, 
    -0.0278448210275673, -0.0822886528365698, -0.0621136149915143, 
    -0.26772553086392, -0.0341516153551491, -0.253197074303223, 
    -0.222765705675088, 0.00429980336495264, -0.242298540989737, 
    -0.186434557070876, 0.106078362179976, -0.220927486575279,
  0.077911805625822, -0.180440078698321, 0.159860596875129, 
    -0.181246608034747, 0.0927758364526124, -0.189854734479849, 
    0.0614386538605847, -0.128460356577877, 0.12191418371295, 
    -0.210299693261295, 0.15799401575717, 0.106553709644251, 
    0.0942017777258605, 0.190305243706267, 0.153064309756106, 
    0.0767846456136216, 0.0986618855187188, 0.16193822927869, 
    0.131213041705565, 0.058296552211307, 0.0814791173348808, 
    0.108419041051561, 0.118383683687479, 0.14317576154569, 
    0.158529184125243, 0.149075418905601, 0.168047233083061, 
    0.206031378288746, 0.172790333285959, 0.125126053548721, 
    0.149956707192913, 0.140832004756583, 0.163382858394992, 0.2684856586461, 
    0.296281113133041, 0.218341868359997, 0.193020346588961, 
    0.293314311441657, 0.282088518435634, 0.197240185186786, 
    0.376374497461576, 0.498816185768035, 0.220451025928901, 
    -0.0771816217400343, 0.215279924272095, 0.618304012826599, 
    0.231061138005841, 0.0353436535316345, -0.0550236460430831, 
    0.274747806448054, 0.371497031109908, 0.436676716251563, 
    0.400239516434093, 0.141558112178074, -0.22951165121794, 
    0.499442627526676, 0.607545702686484, 0.195378708185564, 
    -0.144640477115924, 0.34656164870218, 0.276865101002802, 
    0.370019173780122, 0.447204668379049, -0.0187597108805764, 
    -0.0676551144193317, -0.126015422669944, 0.115704992705599, 
    0.364331611207566, 0.495495456606968, -0.311399733407684, 
    -0.287694866307014, -0.105127706691125, -0.229519158559602, 
    -0.12149944550447, -0.231479515957187, -0.153655034557482, 
    -0.204358351333466, -0.142612970166955, -0.047964728493091, 
    -0.186985496060139, 0.0997996955037643, -0.0856177428395388, 
    0.0811541458025001, -0.0589570358709312, 0.0571167258257308, 
    -0.130070933609127, 0.000317982092860811, 0.0154146643939677, 
    0.131843467896485, -0.112066962679097, 0.165147074512728, 
    0.0197441568499139, 0.00989426261071694, 0.280402319070165, 
    0.205379960551998, 0.0438117706010559, -0.0836690965149093, 
    -0.09001173625323, 0.0929816609503599, 0.396726873082431, 
    0.288384442828093, -0.14323144494994, 0.292879598824331, 
    0.568313775347241, 0.127503476107409, 0.235835562527622, 
    -0.292137305983843, 0.6255104032876, 0.319100161400232, 
    0.151460517748496, -0.16074432525978, 0.571862445474279, 
    0.294728586285135, 0.0724321701971965, -0.154671491742117, 
    0.218599157670635, 0.460557327929596, 0.425496466941032, 
    0.197467432409879, -0.0941542774004191, 0.0959099235741249, 
    0.674059778909781, -0.127876431644298, -0.370245935083952, 
    0.135448014849096, 0.387706358461516, 0.0487063475726606, 
    0.130241692821424, -0.0700940846445717, 0.272902947759585, 
    0.110508032802629, -0.081503747670704, 0.300210702077213, 
    0.479096837926458, -0.0261784439004732, -0.192714433530967, 
    -0.16093890174528, 0.284071740363887, 0.328269254421646, 
    0.0649560934003079, -0.116253140165323, 0.0823877911327342, 
    -0.18923927168056, 0.0163999495607419, -0.119840115124977, 
    -0.00876256989909144, -0.353132421913228, -0.0821785432807534, 
    -0.169272289281085, -0.28672095954013, -0.000273064712368001, 
    0.0657741938472755, 0.113269870397902, 0.128046004795623, 
    0.125462750049075, 0.116819599495313, 0.151661871762066, 
    0.191272317371042, 0.134613327958232, 0.0606740320045137, 
    0.137704703573977, 0.172894970036768, 0.363517727109955, 
    0.397188349716433, 0.181500362816371, -0.0214600263892966, 
    0.400295644455441, 0.530190290319148, 0.184463149802131, 
    -0.144291214328028, 0.274349221526137, 0.316812013588143, 
    0.77778403198884, 0.579335208988209, 0.0393693105412002, 
    0.109187047816001, 0.449840791797813, -0.127159213240007, 
    0.405159548621772, 0.405324582469459, 0.0350680965720471, 
    0.0780681433306365, 5.24268027721209e-06, 0.0411404994235423, 
    -0.0211534905127978, 0.0314423384228766, -0.109743199175449, 
    -0.0263105130267344, 0.0122647969740266, -0.11784328137138, 
    0.0805272857012906, 0.157046038826644, 0.112104496705995, 
    0.0821576422716444, 0.264791726132706, 0.334282432133912, 
    0.229578021767584, 0.169402949448294, 0.174332953448436, 
    0.225475046681138, 0.351690004635159, 0.321164312319082, 0.2642686682804, 
    0.401763393590872, 0.41760894688377, 0.189969426630867, 
    0.124839079010362, 0.576673012543139, 0.31524543737837, 
    -0.0542121810448235, 0.142421223711113, 0.749834598022713, 
    0.29985990676724, 0.514310074462746, 0.406204741968951, 
    -0.422367881683326, 0.221654375803865, 0.417025100314113, 
    0.337132475465054, 0.617051462976647, 0.250420722314961, 
    -0.0141015245055757, -0.121287846565233, 0.125518812069702, 
    0.0626566688099812, 0.0105207870307095, 0.0266048077709305, 
    0.00779827450744847, 0.126073176430275, -0.0461224022204697, 
    -0.0330560141568041, 0.0245120738273536, -0.0269447197863258, 
    0.0546533686119483, -0.0605586836226405, 0.055370162437095, 
    -0.0555246608256501, 0.027291434361832, -0.00935244304423666, 
    -0.0456334598343004, 0.267529727975985, 0.0484783035489363, 
    -0.291971283238182, 0.0839213654984527, 0.522896980045319, 
    0.263163857206584, 0.0842591498878152, 0.00515961205844585, 
    -0.220961982883782, 0.390111620082512, 0.41103353659977, 
    0.143282388488099, -0.000114968534696294, 0.416960506800155, 
    0.180815821410016, -0.0322966982303673, 0.131655479790443, 
    0.322180866006095, 0.013096880749289, -0.0288003281233892, 
    -0.0729667695544458, -0.223158043133803, 0.108682395335943, 
    -0.137752350202205, 0.0711802604309013, -0.153293634290493, 
    0.068138790193335, -0.142168336291879, 0.0744056028755475, 
    -0.230702709483107, 0.0229490038737793, -0.0533070285641522, 
    -0.0256064291240279, -0.0574987553236325, -0.027998671916876, 
    -0.0532427643217923, -0.0519313580625304, 0.058528512920461, 
    0.0597736494664807, -0.295522731479296, -0.217259014335732, 
    0.469709770554007, 0.287176607754606, 0.071750908932702, 
    0.0686354069345634, -0.245764434528413, 0.227042431569423, 
    0.194820349077898, 0.348074163709582, 0.779701170014186, 
    0.296576514070601, -0.0120018991714417, -0.0238337073766359, 
    -0.248508765373521, 0.338037006170322, 0.233323456144833, 
    0.116756287423983, 0.434292608847275, 0.217220092621039, 
    -0.00336046992466148, -0.111157062607527, -0.0820812877987885, 
    -0.0435307121568999, -0.0996260743536049, -0.0671135982860543, 
    -0.053962110960215, -0.0722895260960954, -0.049538232090948, 
    -0.0233520792169281, -0.0494604527983918, 0.209621986925744, 
    0.00396642693305289, -0.11780205754716, 0.0698709032051757, 
    0.671525761151073, 0.369364736709244, 0.143993620094967, 
    -0.237033847593484, 0.31882171365671, 0.229485442816414, 
    0.273204509981998, 0.741440097095039, 0.242679683644506, 
    0.0727114387329114, -0.419148869557516, 0.0109552725870181, 
    0.2232117327096, 0.795456985399496, 0.476483300354892, 
    -0.0324209908798427, -0.159053778598278, 0.104397935938763, 
    -0.24138023737041, -0.0226260067588192, -0.168359869772978, 
    -0.058931997894975, -0.147397011906859, -0.0581190086490543, 
    -0.103943580575569, -0.0668581709829355, 0.0943634237877861, 
    -0.0460319421314508, 0.0920668529771376, 0.166443528545493, 
    0.379315116786935, 0.384848945313327, 0.216486703306161, 
    0.15035577579763, -0.358845332671692, 0.108520732230083, 
    0.503875780191565, 0.405763561094602, 0.213248748033539, 
    -0.300996516734907, 0.0437604422604742, 0.275130533507991, 
    0.778721672991785, 0.59831588242316, 0.140099959282003, 0.113998999343277,
  -0.0369517657484862, 0.0860733666548515, 0.183255993461016, 
    0.183021719621652, 0.140530729580137, 0.113236268612658, 
    0.231900719132895, 0.398706968080655, 0.319099686225307, 
    0.165232248473147, 0.116110112213838, 0.271202902924968, 
    0.566544321059177, 0.45626457823465, 0.184661744479188, 
    0.0286719612574306, 0.631409153750334, 0.639435938049144, 
    0.218965696420752, 0.0240386825191361, 0.617198140726289, 
    0.432321629795295, 0.0360539929614145, 0.248734868198477, 
    0.659781021924137, 0.0609094881522942, -0.163995861766298, 
    0.0710278116371884, 0.480024614103707, 0.146557160234615, 
    0.108412610897286, -0.179017950070008, 0.137179640872634, 
    0.336680222642083, 0.352474782765103, 0.137139946632247, 
    -0.105907083833978, -0.0288986777678018, 0.204258298750453, 
    0.274367381712308, 0.34038680736799, 0.28054214220848, 0.150234111382804, 
    0.103695409247449, -0.0946135784593449, 0.225669530048109, 
    0.432527439908579, -0.0419004526021946, -0.0666370623938548, 
    -0.0707177621755963, -0.0231867496499324, -0.224041543256041, 
    0.177866179446054, -0.132938770696458, 0.0622403538497761, 
    -0.159518472010465, 0.0195771870693049, -0.126654340925592, 
    0.0351679975271863, -0.256902300452029, -0.0166431002777962, 
    0.0424445026212255, 0.0996166821149273, 0.189376890589553, 
    0.208724237424176, 0.147577218124102, 0.129131219090223, 
    0.204631668693621, 0.206074792326534, 0.155020351492197, 
    0.178581811759391, 0.184384314773957, 0.179775106675746, 
    0.212902632797693, 0.222873223613137, 0.149858566674144, 
    0.159891968836976, 0.296839810779929, 0.200681225066111, 
    0.162075259151132, 0.282662130835932, 0.101976250960407, 
    -0.00705656355322075, -0.3026204108294, 0.409538172224634, 
    0.402328743593098, 0.337665578004549, 0.275801007102045, 
    -0.00681674648782266, 0.557404845070979, 0.187378169111525, 
    -0.0999345385940034, 0.263890861932742, 0.261539658270577, 
    -0.169525975019041, -0.0713930321387401, -0.0694675004169706, 
    0.265047182762223, 0.0422158493863991, 0.0148703120923009, 
    -0.0151902805031041, -0.234348624416648, 0.132414556481644, 
    -0.109279966944335, 0.0830325578224503, -0.263688430411731, 
    0.0385242385061559, -0.255220810745356, -0.156040520639124, 
    0.0248132842128556, -0.0731474660513858, 0.280654078069446, 
    0.0595105608448092, 0.207240087901194, 0.322614710367427, 
    0.245359390065955, 0.448334461432689, 0.143128335050626, 
    -0.169978299264621, -0.115198583746885, 0.504112106209169, 
    0.201911213509044, 0.0199861321248744, 0.808954692748996, 
    0.309781047254442, -0.0398738344515052, 0.58155268995946, 
    0.405097272278424, -0.167969111165331, -0.00577910372804216, 
    0.752387694092506, 0.399746859597801, 0.153862557530474, 
    0.105997297832473, 0.0977735107056578, 0.0655921822170735, 
    0.0697253441499466, 0.164693729099942, 0.0706607066235815, 
    -0.03624376865661, -0.0428874606081251, 0.355437362518957, 
    0.140922881825498, -0.0438710770033986, -0.0313101588237824, 
    0.375379593233516, 0.276395262506426, 0.0984215805647465, 
    0.0799995941705909, -0.322214823939461, 0.183441367703393, 
    0.426878415777371, 0.187474140574694, 0.190248902757993, 
    -0.187242008993844, 0.556050283646027, 0.151140348567542, 
    -0.0562017352603222, 0.39874919274066, 0.104614103957243, 
    -0.320235097091968, -0.083773449319676, -0.167615862495666, 
    -0.177348024292214, -0.0885635070815643, -0.205527366747534, 
    -0.0609817729806585, -0.166043249718654, -0.00281318405966072, 
    -0.177553131365036, 0.0826589702669627, 0.00717299051868754, 
    0.0490880533430131, 0.0455395049327965, 0.0618459181853639, 
    0.00473512529147102, 0.0261226074758192, 0.084322285580087, 
    0.105916644469424, -0.0582747626149166, -0.00859707353673491, 
    0.214177734251824, 0.293281284444349, 0.148785150478034, 
    0.0247169885047231, -0.0898641761275184, 0.16581301183846, 
    0.4854675845215, 0.0662374526321671, -0.356279123290489, 
    -0.171871695553843, 0.761663593926243, 0.311331716412851, 
    -0.0354076059642151, 0.0617976152649195, 0.434643102856882, 
    0.82401104046265, 0.445534356527275, 0.116777098150564, 
    0.216185177150339, -0.564255609016568, 0.244044080993955, 
    0.28424735258535, 0.0542227144160744, 0.00909154983414556, 
    -0.0631954860128645, 0.199126441160961, 0.0675060086433309, 
    -0.19690671396101, -0.111240451050157, -0.0956860462742516, 
    -0.137354342799079, -0.0743232326172894, -0.13640766803635, 
    -0.123038454193187, -0.0728436104610182, -0.147507984772842, 
    -0.0681082627940296, -0.133571788541311, -0.0516063499911033, 
    -0.137363505981422, -0.0544854824301388, -0.0266769459074305, 
    0.0273431439917324, -0.120563521921629, 0.0152556354568934, 
    -0.191006018699282, -0.106201311863527, 0.0207267891690009, 
    -0.119520813932551, 0.132376698448563, -0.014509778420462, 
    0.171026440814362, 0.228643481925428, 0.12183286248511, 
    0.0600588309029289, 0.0713061246841396, 0.200646112622483, 
    -0.22245873284732, 0.125669734093945, 0.625867824910984, 
    0.156581454306808, -0.371683363396043, 0.286520746242045, 
    0.544013602458013, 0.140291960063954, 0.0635315982452467, 
    -0.14621887995374, -0.0399460556643551, 0.633469887868226, 
    -0.241477210324744, -0.197828359335932, -0.0821357353741438, 
    0.160017332242834, 0.292109484371473, 0.126560314288793, 
    -0.117868499084578, 0.24270141874138, 0.0745452029964561, 
    -0.228498168449279, -0.0972049568650666, -0.128471913060916, 
    -0.0737693481032495, -0.159266089814215, -0.0564510669471783, 
    -0.181000918406796, -0.0731038223232361, -0.130865336970429, 
    -0.0449225719553587, -0.135636836783993, -0.00215276580104695, 
    0.0664608038848874, 0.0746953952131226, 0.0782155025402036, 
    0.0392960051988936, 0.0558455902669744, 0.0625681831520449, 
    0.0578586486589257, 0.0697252882264305, 0.0246195100101575, 
    0.123978255241025, 0.157576686707265, 0.101580206834574, 
    0.100753655299619, 0.281416738194143, 0.231635712838046, 
    0.122995857114459, 0.102378468434676, -0.140969984209026, 
    0.384782251121815, 0.41415190141285, 0.0936545200765713, 
    0.120651583072021, -0.334066203903266, 0.166007350801643, 
    0.690396921115803, 0.252741863174016, -0.206420263525738, 
    1.03641343019151, 0.494194529217404, 0.0648803298120132, 
    0.054632331223368, 0.0762243578838002, 0.0772583177255079, 
    0.077098686515612, 0.0750326745033145, 0.0733701599759832, 
    0.0879318793628091, 0.0887262335303637, 0.0446810732978262, 
    0.0747102313140464, 0.134752484087934, 0.132055866128359, 
    0.11601150897796, 0.148971376412139, 0.16201194681705, 0.170345034191241, 
    0.210454111449649, 0.194164178622208, 0.164677192591766, 
    0.190355801888319, 0.144117587310547, 0.283453881704254, 
    0.380555478273036, 0.179033009461963, 0.0869908686660534, 
    0.560181663197073, 0.28616132207792, -0.0307736177297581, 
    0.158297035191543, 0.638768544157115, -0.0354128452898991, 
    -0.00052748692824324, -0.337399978088745, 0.225798189530934, 
    0.555722461164103, 0.372893652710567, 0.123561705487685, 
    -0.0255318599010113, -0.0960875659839991, 0.457792996818821, 
    0.0834358748480989, -0.100714643738957, 0.333983957502199, 
    0.0762468924952279, -0.201810649861747, -0.00133616347408067, 
    0.359223162172239, -0.0761140629721674, -0.0709927672770459, 
    -0.0609881262026554, -0.263311591737575, 0.0360322573176953, 
    -0.0852429711718263, 0.0465496869098575, -0.185448842176895, 
    0.0375274104800479, -0.129075033555403, 0.0324635529649616, 
    -0.259450417027289,
  0.27992869772999, 0.245052903823752, 0.21485471532242, 0.278150189967372, 
    0.228187168434019, 0.123205755690581, 0.327573504022059, 
    0.313203117651176, 0.139475751918274, 0.427755835235055, 
    0.366367291228845, 0.0497250498736413, -0.431031486747991, 
    0.456731528355377, 0.630108563250392, 0.0937103416787528, 
    0.0259115820510075, -0.250605397116567, 0.235105480180973, 
    0.350774786114437, 0.212549418287567, 0.27376524250664, 
    0.125806151811739, 0.0317150332156633, -0.0782671008692506, 
    0.115050812661728, -0.104345483679476, -0.134818982134441, 
    -0.11231519057164, -0.115193783188231, -0.162157109771921, 
    -0.242028591178855, 0.0277913052114214, -0.116066850481399, 
    0.017567571674957, -0.1631483306295, -0.0306367464537089, 
    -0.116913685526645, 0.0318734691215138, -0.268694065428064, 
    0.102791612241687, -0.0529457275013964, 0.11349547835117, 
    0.326334521075421, 0.175294245126514, 0.044747050467103, 
    -0.167647612774345, -0.0724899605391681, 0.301224997599923, 
    0.385385301758658, 0.245307647416188, 0.0181792958664032, 
    -0.126296851834718, 0.532247570061622, 0.532579746302667, 
    0.139479209006772, 0.0216084957525799, -0.385956906477235, 
    0.849524029462434, 0.560729249007466, 0.0858662087168429, 
    -0.366483813797979, 0.374372912865557, 0.600964035007943, 
    0.120159323124587, -0.147001348425553, 0.164413247788645, 
    0.40220068486609, 0.329192892407392, 0.206687256012002, 
    -0.155220316930483, 0.315124774745459, 0.350623569550928, 
    0.071443890031516, -0.0553403224005994, -0.141620964488422, 
    0.440444170772713, 0.19481421223396, 0.0237143434887871, 
    0.0197236358378066, 0.172197223764765, 0.23620208516231, 
    0.160732723294549, 0.0870571088495826, 0.029237312013037, 
    0.0648892130370944, 0.246844254618848, -0.0469356868489394, 
    -0.131668276183859, -0.149883164076373, 0.175628108386753, 
    -0.1737452710249, 0.142305699730481, -0.128694206826921, 
    0.0885443442286277, -0.1038226921654, 0.108098012001813, 
    -0.167774593137455, 0.0897536780400027, -0.115219129292965, 
    0.166857619145979, -0.0302072745747619, 0.0384296334749206, 
    0.0193606344151729, 0.058339686748531, 0.0351251540209698, 
    0.0708461500204394, 0.0289042650637359, 0.0253847436787812, 
    -0.10245202457911, -0.0111030759304292, -0.051478299179352, 
    -0.0462691790411361, -0.0314442837173451, -0.0365905712993227, 
    0.00539218300570595, -0.0454899908717927, 0.0394290462534056, 
    -0.0377164022964479, 0.0050613544030328, 0.219215380606136, 
    0.0672012920175482, -0.205090782593881, 0.0718682774814844, 
    0.37940966897505, 0.274291233764329, 0.505386094278658, 
    0.287374115343223, -0.419652339084352, 0.119711145063526, 
    0.508237827396722, 0.0963389808489499, 0.499350108241383, 
    0.628725482494571, 0.283052809156702, 0.216659732583611, 
    0.383591561627686, 0.375447723349484, 0.239701050038226, 
    -0.0489903250098377, 0.269988638285387, 0.209187430916822, 
    -0.203281397980306, -0.159013116209803, -0.0803963665074457, 
    -0.181886240305011, -0.0435233086972986, -0.145290502879994, 
    0.0221742305912914, -0.176990746160583, 0.223939312513899, 
    0.0861595782123802, -0.00834148883894613, 0.322894244103459, 
    0.317416033770292, 0.123301168730218, 0.0616478965416793, 
    0.389459475127113, 0.313239919985524, 0.122970624575568, 
    -0.101416557053492, 0.540892596789855, 0.277046274291643, 
    0.00861449181320963, 0.321468539685323, 0.377473353751372, 
    0.0250610622206572, -0.013066993766873, 0.595456704928876, 
    0.261297894432178, 0.0252439331425593, 0.0321758873763347, 
    0.00821862464065368, 0.0198346193255432, 0.00987668604972663, 
    0.0174353918956386, 0.0139566008160772, 0.0168842939652002, 
    0.0216638345713484, -0.0118467285770105, 0.0634943331370547, 
    0.0844684539864468, 0.111987961676673, 0.165930958798241, 
    0.183930015721094, 0.157220228396645, 0.1495908857375, 0.17868321413968, 
    0.156209644209845, 0.118282864836855, 0.206564588136231, 
    0.219009562048573, 0.142926647914804, 0.19886718405223, 
    0.358028624416068, 0.249586927325361, 0.116583030032076, 
    0.302173962857779, 0.390973707522962, 0.163822692101463, 
    -0.083113236818839, 0.381452715620117, 0.539975845926184, 
    0.0432089600718718, -0.0450881129765762, -0.189311872609309, 
    0.579306350285535, 0.24152223033061, 0.335613012523742, 
    0.353733652263283, -0.255005815196394, 0.302488895274942, 
    0.314697248814968, -0.0301784687507918, -0.0448682296299862, 
    -0.20332679532002, 0.620891291413591, 0.195679851269063, 
    0.147345336327453, 0.218319023525869, -0.121756250618142, 
    0.1856780935938, -0.233110726307548, 0.0916796206161232, 
    -0.417710692144475, -0.160843461911151, -0.00877210321158978, 
    -0.138876271442772, 0.224527177773064, -0.251882061753749, 
    0.0459491381883684, 0.117518975173466, 0.141601844386406, 
    0.0755100385861248, 0.0771720661604528, 0.101983582050162, 
    0.0958289963999506, 0.0919726469352456, 0.0801660685526418, 
    0.0121184269701023, 0.0333435591584384, 0.0604500539958286, 
    0.064280056960855, 0.0653046445566151, 0.0704903049925117, 
    0.068806479949089, 0.0690722342012103, 0.0987284406180354, 
    0.0806231054691105, -0.114888910936212, 0.329545521480494, 
    0.251070358586378, -0.0676013675600199, -0.198698952912654, 
    0.465348183683975, 0.537817423570841, 0.171037632671835, 
    -0.103441244625057, -0.160089837448508, -0.397343105999129, 
    -0.0837233774618855, 0.709792240702648, 0.168484560628803, 
    -0.0683108757294574, 0.464058776496518, 0.281880997071902, 
    -0.547909124440614, -0.502704562425455, 0.0575098159325745, 
    0.524647855317592, -0.210639730748336, 0.0105653527015689, 
    -0.201324468592895, -0.0650324430949773, -0.163067434338095, 
    -0.0898268622623783, -0.147305798866249, -0.0776136749236481, 
    -0.100720733978814, -0.14391477698966, 0.0533434802747746, 
    0.203153857811023, 0.232177641556568, 0.0130016271367018, 
    0.00330246044685041, 0.452629808210043, 0.483660747819302, 
    0.201179444244933, -0.267729192638513, 0.252171670628508, 
    0.554326138184249, 0.144713834927183, -0.282866111608818, 
    0.124777761217489, 0.631460489790654, 0.240331561157741, 
    0.0750957553236701, -0.0918390053741397, 0.317213977790091, 
    0.263805790230914, 0.305252507617371, 0.695833178386875, 
    0.389799239969407, 0.0832060635606215, -0.267543110117795, 
    0.15438160878035, 0.472760610553004, 0.152671808194056, 
    0.318948571722435, 0.616308256683697, 0.0292510575373648, 
    -0.0550126364668346, 0.0353429639029314, 0.432066793928262, 
    0.0260818041008752, 0.352724081929065, 0.570554545007959, 
    0.139621530091053, 0.0815233019248737, -0.030693482088914, 
    0.246795599872288, 0.201838171004713, -0.00384109035392004, 
    -0.0290528677658708, 0.076005414591585, -0.239462811906603, 
    -0.168118885140539, 0.301445318429914, 0.24163230398325, 
    0.0248900197840377, -0.129653653924259, 0.123083507202836, 
    -0.430561197771327, -0.151891598867182, 0.0144591412379341, 
    -0.201617976258741, 0.128708901799375, -0.101670607498579, 
    0.110509649743004, -0.245547224396824, -0.000163553761937801, 
    0.0918483127563978, 0.149552423768171, 0.129455063172547, 
    0.128585683323118, 0.289876797928232, 0.340676065304991, 
    0.224169714084449, 0.137345243893773, 0.176817010987645, 
    0.311212435389834, 0.333711630731301, 0.29655630621368, 0.28912076923353, 
    0.293242601224568, 0.257768237419139, 0.22418216851909, 
    0.248180343984138, 0.277053418601372, 0.281122727226867,
  0.771142064321767, 0.344246075505045, 0.328548362861347, 0.200194895296714, 
    -0.323265269568207, -0.0830775181446554, 0.633026896370247, 
    0.200220791469334, 0.24653566819773, 0.92182140197364, 0.285290748435384, 
    -0.0433288423553949, -0.0689264636294254, -0.0881966131243885, 
    0.302265703652816, -0.067151645941394, -0.230098779390148, 
    0.141689558779674, 0.0291238302609434, -0.16808709624641, 
    -0.10735262569498, -0.120491605560857, -0.0788430790965761, 
    -0.115479848695583, -0.09610083240173, -0.153659437761206, 
    -0.139308590024975, -0.0778434770223118, -0.179713577848602, 
    -0.0827690154835885, -0.20045234864826, -0.0559381535666668, 
    -0.0864964486039186, -0.102868769025669, 0.159373774779742, 
    -0.179944619535155, 0.0615486257699361, -0.128515140328053, 
    -0.00887385178160541, -0.167717689786068, -0.0655940404007244, 
    0.0952394711389467, 0.11529737925109, 0.0678981112765362, 
    0.0940399510236869, 0.156347636900668, 0.208404498765787, 
    0.242329991327135, 0.165259282331557, 0.0562710730314155, 
    0.149509636662986, 0.238846760684719, 0.17817356455275, 
    0.408179948690635, 0.559394224752712, 0.244314530900467, 
    0.0364727939800634, 0.615660259063677, 0.36104762321122, 
    -0.0385504287876845, 0.360807589845835, 0.56552258953605, 
    0.475912734734098, 0.298210198053904, -0.187125344041551, 
    0.318004997106066, 0.531713119367922, 0.23306344703984, 
    -0.0491786683576186, 0.317894154438785, 0.29775606470188, 
    0.156166247493965, 0.112761784172362, 0.0815838505009947, 
    -0.131284850543417, 0.190563685755918, 0.0761500730379282, 
    -0.0580120705349779, 0.0864028712439194, 0.158379308349886, 
    0.0247955792153229, 0.0125169030733271, 0.0113115320405742, 
    0.0139476839356677, 0.0149218509327676, 0.013191905008577, 
    0.0145373527784314, 0.0205078388341537, 0.0224236182881208, 
    -0.02375489511829, 0.0494021529711983, 0.0458290600531442, 
    0.206101724929086, 0.229063330204717, 0.101231545280131, 
    0.0662424447404108, 0.251652776794369, 0.260880119890897, 
    0.26819912321828, 0.105047565288335, -0.0492082278238319, 
    -0.0251748967238224, 0.259939419122777, -0.0125444110991928, 
    1.01542187425179, 0.445594326030925, -0.199363037152338, 
    0.433174520012282, 0.821760975937446, -0.221170122429949, 
    -0.129413879466479, -0.0585183909145566, -0.11243258851238, 
    -0.023373721985211, 0.0033348090878238, -0.0528812611084327, 
    0.009051815873695, -0.0796690471506556, -0.0599715289174532, 
    0.00135210540140152, -0.123008365636072, -0.000984159361188591, 
    -0.0963538274281962, -0.125486290952116, 0.0789925221720186, 
    -0.0364253691065295, 0.050664918944473, -0.150821370398701, 
    -0.0117935959833013, -0.046700580938085, -0.0102560980291079, 
    0.00402801198892937, 0.137439606104343, 0.0546980858648513, 
    -0.0132870689811337, -0.000201997125896483, -0.00310850768568396, 
    0.385757405264538, 0.0754239705419964, -0.371925408247508, 
    -0.053383985286584, 0.58858701195794, 0.135941675596793, 
    -0.0841221817772892, 0.205151568427875, 0.554165444403417, 
    0.28546526653406, 0.411268011641268, 0.991051252827485, 
    0.0548204096263808, -0.375166231343945, -0.157197861849811, 
    -0.120206244504002, -0.194021418301457, -0.0224239623500622, 
    -0.174694404024849, 0.0762535773082942, -0.237650395728551, 
    0.0386343965002346, -0.11683617608742, 0.103979105119345, 
    -0.0432548453377472, 0.0724174207150467, -0.0522270785414613, 
    0.0748072954136601, -0.104574242562821, 0.0374016603733943, 
    -0.00332907401108623, 0.0469022880163936, -0.247959374309448, 
    -0.0114521040272768, -0.087036898685578, -0.0805322693605496, 
    -0.0580626831131138, -0.058371473088477, -0.0810809558708133, 
    -0.0715822039458109, -0.0640464332258382, -0.086301908925683, 
    0.119845133462039, 0.240096322171708, -0.0769587201081097, 
    -0.0675338368525631, 0.714127952496271, 0.30442987519371, 
    0.380057805215305, -0.22844223699386, 0.696415602828719, 
    0.275055956646858, 0.0661003617804569, -0.0866748833113139, 
    0.249974291952144, 0.118429354090208, 0.382070035917652, 
    0.801678374661914, 0.278606580833197, 0.0888866351041858, 
    0.475256426928694, -0.0078707013215856, -0.164003850751196, 
    0.136190573434648, -0.0968911568908152, 0.248723239644485, 
    -0.183690189374714, 0.192576805425608, -0.512193756973915, 
    0.0173966127673009, -0.313787895960986, -0.0626327469901144, 
    -0.274615501531831, 0.0281319005623039, 0.0933345052754582, 
    0.18317838846581, 0.246601196756749, 0.203384658360863, 
    0.145985803327179, 0.128616018404186, 0.237210921678771, 
    0.332323661748275, 0.171036612012917, -0.00383723519916771, 
    0.0417903773155543, 0.128630045609467, -0.157001369013946, 
    0.0821417493665001, -0.0962008286465869, 0.0040460236828293, 
    -0.061225543378821, 0.0509993415633437, -0.119367367087743, 
    0.0221099217643935, 0.0496482492495082, 0.0707815808025934, 
    0.140214945758714, 0.165045999411882, 0.112177233330546, 
    0.0825202067764799, 0.167777686234681, 0.174642097413517, 
    0.134775183765943, 0.150181962828072, -0.0287194358516584, 
    0.117793876684089, 0.542422756971248, 0.28779978883288, 
    -0.00380743804323244, 0.30195297823412, 0.670488315137091, 
    -0.212705510183359, -0.068783911836317, -0.285968628806208, 
    0.143274955241295, 0.766431574933967, 0.0666968539734828, 
    -0.292972790755674, -0.124925365835968, 0.627447590488296, 
    0.218535677405691, 0.0821888267037912, 0.402075382219222, 
    0.187014997495335, -0.243921205297758, -0.131837726949317, 
    -0.0115732721418864, 0.22779470316419, -0.0964016354833958, 
    -0.0640438951106266, -0.13704766371763, 0.26603616101736, 
    0.0747614057765177, 0.000237486972986423, -0.0291183921608541, 
    -0.00661647989701424, 0.113200046736748, 0.104580747328537, 
    0.0658966861005238, 0.0932258517522392, 0.102665958096746, 
    0.0216977332287402, 0.061194158246936, 0.341146980691506, 
    -0.189189771007433, 0.171148893016817, 0.508116230462047, 
    0.192847636671448, 0.0619309554666379, -0.00435946088364005, 
    -0.261763986832506, 0.29230742281174, 0.448219493499697, 
    0.239598894208639, 0.163795692034536, 0.153549759621279, 
    -0.183627445033378, 0.487621635383999, 0.0890947525458362, 
    -0.123970277850785, 0.241659790050652, 0.241820552105568, 
    -0.0164139396351092, -0.0633372063232928, -0.209145569814794, 
    0.0667626496709239, -0.109830504598046, 0.0395250710333289, 
    -0.124933171486934, 0.0500711999409282, -0.143382265944957, 
    0.0344463480998143, -0.211923339371598, -0.0342543435166704, 
    0.0974071701332151, 0.0687037576281201, 0.126334605037486, 
    0.204844306270312, 0.0692301906758672, 0.16036893254576, 
    0.32349703870905, 0.147731807692897, 0.26161268594892, 0.249365551583813, 
    -0.0585456384119508, -0.224137022863899, 0.629903706300479, 
    0.237357979099847, 0.00964617248413864, 0.0336315541756208, 
    0.102963269177596, 0.358952164031885, 0.685742680952967, 
    0.26380858450297, -0.00512852038784176, -0.0635673590285826, 
    0.0304247970449179, 0.142600657324788, 0.0126486828049957, 
    0.0585271995607508, 0.196786128570704, -0.100000040232255, 
    -0.0427237586139135, -0.218878716345349, -0.0936432506581529, 
    0.00227286957534324, -0.141017916897076, 0.0555832409577449, 
    -0.0161968613674329, 0.0596014487479152, -0.0286785373585735, 
    0.131302357656117, -0.176689569251806, 0.0838471638852451, 
    0.123117882793929, -0.00149671079881068, -0.039239501362154, 
    0.300386457057738, 0.167853518891107, 0.132680065962761, 
    0.164478850218886, 0.00137229552465956, -0.217449074249404,
  0.35154108763419, 0.0424573607935092, -0.0700433143413918, 
    -0.0946373423293234, -0.00542734418545342, 0.0636871760809167, 
    -0.0234453619938372, 0.076827437490903, 0.0369057116186486, 
    -0.0537932458772126, -0.00787934682068479, -0.0635930167702583, 
    0.0135866702644101, -0.0291804628610954, -0.00415132717960629, 
    -0.0573162819982547, -0.0201408725949737, -0.0057784616295859, 
    0.0529434712602136, -0.11197478481197, 0.143589853201547, 
    0.351375138724182, 0.282260251790522, -0.112673526513314, 
    0.328375003724123, 0.328943194440815, 0.0895024302900769, 
    0.546911895023137, 0.248846465594972, -0.194926231010202, 
    -0.54703961388231, 0.142279303296382, 0.928486652652141, 
    0.23277218541087, -0.0732881562724582, -0.0947170627981715, 
    0.591444632562705, 0.248515755771413, 0.118013890603858, 
    0.912140060331486, 0.377021220942875, 0.0884511764008087, 
    0.0324934747271737, 0.0484020287693624, 0.0947845969631869, 
    0.0774034578071235, 0.0584872402761834, 0.0780455225984034, 
    0.162484263253264, 0.116944005284416, 0.0581466488153458, 
    -0.00733899053170632, 0.357570622333994, 0.224214386436462, 
    0.0856261050561498, 0.443984182981, 0.332773870760042, 0.124756625314299, 
    0.164347586075562, -0.383309375052923, 0.329341138208437, 
    0.470919276685702, 0.183999240393626, -0.0946845121469287, 
    0.454738423333669, 0.232474970078445, -0.0212943981191486, 
    0.194091079158971, 0.425199912311869, 0.0245059628612869, 
    -0.0657192281643298, -0.0924667335700893, 0.0240851089186085, 
    -0.0331753918869702, 0.0170449805088162, -0.0764098670253398, 
    0.000388048389529619, -0.0304839657159927, 0.0156967998795034, 
    -0.0937712208362087, 0.0148473125496244, 0.0286762849036515, 
    0.188446617045523, 0.259931361791138, 0.286299303306111, 
    0.230051061982219, -0.159938099574241, 0.560035393308605, 
    0.168302890781295, -0.213701118874103, -0.206951613594185, 
    0.58562967388001, 0.664826688810069, 0.214521371517763, 
    -0.18711168107396, 0.228356374156432, 0.00448630406704306, 
    1.04724544308218, 0.332316828546735, -0.337318025573849, 
    -0.259594358559586, -0.0552569600970923, -0.00826930763696416, 
    -0.0119369604319983, 0.0452008492123149, -0.16809980970924, 
    0.107977787128243, 0.377743301984913, 0.0464188539578778, 
    0.0240886520833289, 0.00101134993911295, -0.267935559195193, 
    -0.00285927789564837, 0.0908916063763832, 0.214267245885526, 
    -0.0481493000315669, 0.298543137203834, -0.513703476993354, 
    0.0591526698938788, -0.292716411581186, -0.0835871956157873, 
    0.0490037844865395, 0.0971794322835048, 0.11711784201976, 
    0.111796133885483, 0.122513329319414, 0.112747261653848, 
    0.0877007641919356, 0.00271556885776719, 0.0699660564733882, 
    0.363721166077847, 0.176277197754615, 0.0332656012934683, 
    -0.106368589956625, 0.423825313692307, 0.339965116436127, 
    0.225232727815827, 0.430190508993264, 0.245553778198703, 
    0.392385427295312, 0.70464812698312, -0.0368580753522294, 
    -0.350741563645258, -0.164812200587172, 0.596270953511351, 
    0.194252044939567, -0.00470184290508637, 0.105228250262775, 
    0.715206178354488, 0.0167160722776072, -0.0787944771414717, 
    -0.0862480407643268, 0.129345485334429, -0.239208586228647, 
    0.0403654977935308, -0.33448133701915, -0.132852516290526, 
    -0.140812718069484, -0.135039549328641, -0.176681343955127, 
    0.00188956426724334, 0.107023976725508, 0.166114052485016, 
    0.193903153319289, 0.263931268431245, 0.270147862117435, 
    0.194400745042654, 0.144417768409898, 0.220843080039628, 
    0.314350150493022, 0.296192602151219, 0.243957002310429, 
    0.218958779208483, 0.226721524583699, 0.219535373678778, 
    0.175676677983095, 0.200181326528089, 0.300187024620683, 
    0.207549161491371, 0.0443598958138376, 0.0465386049854657, 
    0.403842910374057, 0.313240453603299, 0.111027599864548, 
    0.00121739033084539, 0.387777402109627, 0.259415807516317, 
    0.0771336084774821, 0.535041878984858, 0.385014836814801, 
    0.18833718128666, 0.252799459928333, -0.16171742465439, 
    0.652173432798328, 0.37794983072168, 0.547830140293973, 
    0.416614094515957, -0.117429161868803, 0.465172729592176, 
    0.233559416720064, -0.332481061920994, -0.0244910222132275, 
    -0.217078621835115, -0.120137180688862, -0.176580236287695, 
    -0.139508995881147, -0.15410140775342, -0.0715014842395627, 
    -0.249931279446909, -0.0382912600651872, -0.0134254090457276, 
    0.0965353692710376, -0.0544799236455655, 0.0332100455551373, 
    -0.0317964247449299, -0.0227512346527099, 0.0484190404272835, 
    0.0112637604258723, 0.0948957572342291, -0.0393705482786637, 
    0.0326285784007362, 0.110743056619441, 0.201014248802521, 
    0.156655688401322, 0.0628139450130237, 0.101371892625407, 
    0.293001447854778, 0.28248073764236, 0.165964542754486, 
    0.116502679512871, 0.238998426578437, 0.249718468113389, 
    0.15596347179914, 0.293846550083064, 0.479591841414926, 0.26260409784714, 
    0.0327550363216116, 0.307218226539544, 0.500440475305011, 
    0.126951612755642, -0.0274226778347781, -0.0670895529020276, 
    0.57436323145016, 0.206426627653364, -0.077645570410893, 
    0.168966337357946, 0.454253683220732, 0.185977749142601, 
    0.0536121880667126, 0.34240263678011, 0.293893536472459, 
    0.449592346777209, 0.411317858663698, -0.149183100791627, 
    0.192197948896872, 0.977343599820159, 0.0597100765627158, 
    0.0104220830978955, 0.430333094678591, -0.124258151568916, 
    -0.311734464986038, -0.0173542483877315, -0.224776891686354, 
    -0.115000242011446, -0.180453491730888, -0.167615509178956, 
    -0.0213226830200836, -0.200382780823353, 0.08762435816309, 
    -0.182116918172135, 0.0822249356266532, 0.0163031941972525, 
    0.0675431755042066, 0.0137984928292818, 0.0453040073142916, 
    -0.0207706979716106, 0.0164905842314403, 0.0271974792861663, 
    0.00956585577030104, 0.0184270605280846, 0.107653015193891, 
    0.116149961107181, -0.0321507749182219, 0.183686446341027, 
    0.326331683562313, 0.137955325672971, 0.0620081820833647, 
    -0.0950124473729898, 0.0646994371138148, 0.101301036682081, 
    0.617015654073038, 0.509623237692002, -0.335292389161167, 
    0.641965265995313, 0.681313449326713, 0.357895258931574, 
    0.295042754718976, -0.0647138001067593, 0.527761743137058, 
    1.07849749361725, -0.0671764455402631, -0.136151844865466, 
    -0.101588916790883, -0.0935140673937674, -0.114705185539733, 
    -0.0323206310574405, -0.00914802045261799, -0.0828378251099024, 
    -0.167136453154111, -0.151461622325028, -0.0388690896778603, 
    -0.0802446072026941, -0.0742597988148964, -0.023029158393139, 
    -0.0904362046868513, 0.0382962887355028, -0.099214451562394, 
    0.0711599414310561, -0.0956867824536228, 0.0350163575102812, 
    -0.0294934481367467, 0.0272453835476265, -0.0137721144035644, 
    -0.00897031696577953, 0.0216241684871325, -0.00929725520760354, 
    0.0221037334205697, 0.0137614073475691, 0.0571474794373147, 
    -0.0217637343547962, 0.0615354193674591, 0.101497701105894, 
    0.093188390643518, 0.111943013629939, 0.128367992979989, 
    0.101373165773249, 0.101520162348636, 0.143184150214209, 
    0.124010645850279, 0.0796581707447565, 0.140588093720211, 
    0.15222018516362, 0.136172973652475, 0.207951802190114, 
    0.326887300094321, 0.292210385251901, 0.153243749533883, 
    0.0154020181715797, -0.000699316190665753, 0.574810756139337, 
    0.304016154737065, 0.0691399818082581, -0.281011034474735, 
    0.190329684217032, 0.557556982088936, 0.317433477461343, 
    0.128232291706022, 0.0707211758458242, -0.244428790136654, 
    0.320048091231318,
  -0.0455210618563821, 0.668725732096309, 0.279676608739737, 
    0.137401812501985, -0.277618381459763, 0.416394268824566, 
    0.323921849023582, 0.214698506937525, 0.601653292301987, 
    -0.0369247616469252, -0.420743758402889, -0.224334023644799, 
    -0.0446074907417118, -0.377697141517936, -0.168026321998858, 
    -0.202944009344384, -0.149802683312385, -0.195100774947302, 
    -0.170937333648158, -0.118207688696625, -0.304754237890326, 
    0.053718407774344, -0.023920176427309, 0.114840651031072, 
    -0.353044381972546, 0.112165984955, -0.275371054962881, 
    -0.0713080766571821, 0.0647960250487236, -0.609858720031087, 
    -0.197559109851043, 0.0322972563963867, 0.0367844879677303, 
    -0.0090464643177355, -0.0987341729288021, 0.0431906735207829, 
    0.170349136438745, 0.129799422342763, 0.0593834408765947, 
    -0.0150766180858211, 0.07119321486589, 0.082550430756627, 
    0.455939283669628, 0.375437421065733, 0.0160338521014569, 
    0.240241174504183, 0.83976534533893, 0.245569050884387, 
    -0.173784372043997, 0.388888479869898, 0.530126004173395, 
    0.156488722247454, 0.0815586204984634, -0.0520497231547621, 
    -0.20724130605319, 0.595519932653549, 0.180856617816067, 
    -0.0624560990077289, -0.0461260565910326, 0.474868975382524, 
    0.241502587405054, 0.0334470801999484, -0.189707850425626, 
    0.0679150898272024, 0.19760164370652, -0.0970382324381967, 
    -0.0938948361417886, -0.0870921359617264, 0.164500201311276, 
    -0.00607232203520007, -0.088730773081709, 0.0397994054759069, 
    -0.054192067586379, -0.00961643544952053, -0.297782741978978, 
    -0.028355420346897, -0.0684560623537002, -0.148564935001302, 
    0.116584425938372, -0.20545543897289, -0.0163138730215036, 
    0.0498238623478352, 0.235919249348875, 0.213048063344681, 
    0.0807314260997219, -0.0022408561287113, 0.287093753893904, 
    0.398138692914123, 0.21974723466678, 0.0914229844278096, 
    0.148924905457827, 0.328843012683559, 0.355656844173926, 
    0.300810369205432, 0.368122115873819, 0.462104615988307, 
    0.37678039403477, 0.240069895473328, 0.232182558778643, 
    0.406248431129699, 0.406958845039976, 0.239562568868703, 
    0.176609022805645, 0.438289148234339, 0.409949141113736, 
    0.150675394504681, 0.0864865561772679, 0.513954029688866, 
    0.266687004796228, 0.0640846155639875, 0.429625171577739, 
    0.44778120852747, -0.355936381051425, 0.501067202938366, 
    0.401135702893752, -0.0119039624515684, 0.0358056357904182, 
    0.600168390456849, 0.510320243622787, 0.173553177073787, 
    -0.139807076488573, 0.0653270002857176, 0.145768442814785, 
    0.531825345239267, 0.137882559471887, -0.166476646206589, 
    -0.223118124169745, 0.0168187772072239, 0.278796028798415, 
    -0.105385116219574, -0.0505490933541855, -0.0253121195347292, 
    -0.0529765500388117, -0.0335523953291318, -0.047261832391889, 
    -0.027233438876081, -0.0452243583009214, -0.00461796231985198, 
    0.141105567674262, -0.186936619779027, 0.458012343663711, 
    0.140798177302184, -0.137565187775811, 0.141146425304119, 
    0.239274530263322, 0.245022405878428, 0.65942254134749, 
    0.216874437646382, -0.067499407760943, 0.0423381729978886, 
    -0.0609102200157697, -0.217229882972043, 0.20191275810099, 
    0.230688197779979, 0.312370805685874, 1.03843463949892, 0.47092783447942, 
    -0.0263252435253852, 0.485335801046134, 0.458050266160124, 
    -0.0866213873644809, -0.0523979025920788, -0.0205835568772686, 
    0.149239293749563, 0.127858921807331, 0.0526290520807029, 
    0.00573108699434251, 0.175685339867832, 0.125566486946586, 
    -0.201060750328932, 0.113287096405771, 0.375971358786866, 
    0.0887817755600683, -0.132688550265922, 0.0464697379283745, 
    0.421362000229328, 0.308490404817872, 0.134052283720873, 
    0.0352754058951938, 0.513779183431628, 0.131623791404601, 
    -0.0516689674448327, 0.0019658235108944, 0.327853609557861, 
    0.202665472236732, 0.0695353001260926, -0.0839603294793522, 
    0.0918963903501226, 0.17159540097681, -0.0772396303135301, 
    -0.0802217206055885, -0.118224736341784, 0.115771527252647, 
    -0.123131171555911, 0.0917563028278446, -0.233549283451145, 
    0.00458053842270416, -0.150549574572252, -3.66879784094443e-06, 
    -0.243532601156524, -0.0594343194104351, 0.0656367183176166, 
    0.0969384592980759, 0.0916951540533082, 0.139064134060708, 
    0.112399685954332, 0.0495681583758104, 0.253384916587978, 
    0.257650550505659, 0.054945208451291, 0.105164661665883, 
    -0.250154226676544, 0.439353294070998, 0.459230901235751, 
    0.0913352551487078, -0.121765567256182, -0.158484042021218, 
    0.560635096774868, 0.22953876562673, 0.0797124406743781, 
    0.0261359514424803, 0.0619482461820697, -0.13901146305733, 
    0.837001614892844, 0.219404573118273, -0.100325471792713, 
    0.0554522387159307, 0.590202723092123, 0.211186799404148, 
    0.0118073418771432, 0.0959659379391982, 0.280434754449564, 
    0.11800265942319, 0.0493421893637495, -0.0412311493948451, 
    -0.172721958329561, -0.106445840986717, 0.0293626197855961, 
    0.178741654817957, -0.14509894239769, -0.189376089806168, 
    -0.105354105741577, -0.123572801770686, -0.13875176608858, 
    -0.104753375637395, -0.143143403047689, -0.0740363080731658, 
    -0.134623797277463, -0.0065142834669895, -0.158253761278647, 
    -0.0062293887018523, 0.0598514728569626, 0.0827856780324039, 
    0.112102164493119, 0.134404786869117, 0.108894099345534, 
    0.12261522822002, 0.173236725895702, 0.128334339204138, 
    0.139828709567981, -0.227715360518583, 0.5267953867741, 
    0.380850543885743, 0.0748375402462659, 0.0141146531619095, 
    -0.268923186967326, -0.0129877524864184, 0.780703749118353, 
    0.223296246985194, -0.170239382591621, 0.113004261276853, 
    0.651840009061919, 0.289146668205428, -0.0552038416338129, 
    0.504418925666701, 0.797541241652235, 0.214989138746639, 
    -0.271444517522388, 0.222670142878403, 0.514515993505444, 
    0.130922967205792, 0.0567195656774223, -0.0820417579558255, 
    -0.0193877554890893, 0.281316966210719, 0.161561736885771, 
    0.0996507984106255, 0.24077729605866, 0.175795436575051, 
    0.176880019231715, 0.28771802584436, 0.123533501437704, 
    -0.118498598060214, 0.607516776976477, 0.310225180770554, 
    -0.00189987159448929, -0.114980826347707, -0.0653494839668758, 
    -0.155983174887654, 0.577738214382971, 0.28621465305684, 
    -0.0974832683899226, -0.0363196642945431, -0.398589472927528, 
    0.204301617947773, 0.469945670479228, 0.223336538761218, 
    -0.0483405413625142, -0.204088692897168, -0.13097585779878, 
    -0.0657709838173488, -0.357878830409664, 0.0717604796538137, 
    -0.325655299782983, 0.0691455181745009, -0.265916923541249, 
    0.0955666981981505, -0.188927330093815, 0.124207522765142, 
    -0.284638919338661, -0.0111763683845291, 0.0875113569355552, 
    0.141321218777308, 0.230720318398828, 0.258845100609633, 
    0.163898242456757, 0.117458468692198, 0.314573154603367, 
    0.356818331333027, 0.181269709618246, 0.0461043051848015, 
    0.0230430041415712, 0.0466978040621793, 0.0603450558500588, 
    0.0912666556540433, 0.0435142891118001, 0.0715354768058383, 
    0.103134358472126, 0.0911987315929179, 0.0213507085037774, 
    0.0503043629472699, 0.0733031509762871, 0.078843556148674, 
    0.0771946847921163, 0.0832274723005834, 0.0713361466864998, 
    0.0686594897833067, 0.0993617151493118, 0.0919086690811817, 
    0.0278468536598151, 0.0576645853258573, 0.135539275186127, 
    0.2674389899632, 0.211234509671252, 0.0623706580900858, 
    0.0775986097034282, 0.437542418179682, 0.203198522255289, 
    0.0126573412371157, -0.167178776089336,
  -0.194505416190631, 0.0566775945319974, -0.374457813116822, 
    -0.113739120607899, -0.167080858718634, -0.245307220135158, 
    0.0251920126119114, -0.302496382174655, -0.0237554054531844, 
    -0.210878696742427, -0.0671312001095736, 0.0774595545502246, 
    -0.058618869703866, 0.0219517970389059, -0.00653994721924762, 
    0.0136020488767386, -0.0750794291742679, -0.0213232225376437, 
    -0.0326470969923791, -0.0933620314708881, 0.0241618549250895, 
    0.110458543610893, 0.0856356179457003, 0.0841285312258885, 
    0.154909882090056, 0.122919949746273, 0.0759110191719427, 
    0.227036455567576, 0.238676971238737, 0.136282178600557, 
    0.155582125700585, -0.26761523295367, 0.223061649781575, 
    0.494851856203744, 0.0623745085348597, 0.0782136415886878, 
    -0.274970961276018, 0.39405697289688, 0.360768667138414, 
    0.126352197753587, -0.047893948335751, -0.124853612801916, 
    -0.147468654996586, 0.532271277048181, 0.371285843346411, 
    0.084630138939819, -0.23591864458955, 0.0278898527246108, 
    0.420845748594582, 0.227596043553195, 0.0943940970580293, 
    0.214707680551766, -0.0104941200355806, -0.0339961004218759, 
    -0.0106168834900018, -0.0949272480549539, -0.0458350341768063, 
    0.135701176114367, -0.128469544955174, -0.073399721281071, 
    -0.121951798755525, -0.0718330202612044, 0.0455441499216038, 
    -0.221971909511293, -0.00841435199552498, -0.363608324859085, 
    -0.191753400064488, -0.0329580201956302, -0.217620861018337, 
    -0.119211746735268, -0.0270832052604928, 0.0602468526889776, 
    0.0855587601691777, 0.091414945010851, 0.117751939259013, 
    0.117050985951688, 0.142525645747119, 0.172383601306183, 
    0.0950842035278742, -0.0144048919780725, 0.129062955291524, 
    0.26887719764701, 0.20395756490417, 0.14041062006701, 0.132638638544391, 
    0.347515332176636, 0.537553171641288, 0.225693885342068, 
    -0.167718851745818, 0.242754392767854, 0.534635075074561, 
    0.365321492816173, 0.201095513199141, -0.309821862959432, 
    0.106155871604691, 0.483803519378546, 0.103300408467509, 
    0.0341698563585392, 0.0916097446015122, 0.526685795431776, 
    -0.161044640799005, -0.104201886154104, -0.167186634095853, 
    -0.147616951241655, -0.164636896891062, -0.13298892103796, 
    -0.171553098370628, -0.119695318775032, -0.129126916576196, 
    -0.124833833645034, 0.0376823850576678, 0.0324169620065985, 
    -0.0301448797503876, 0.00773750719062359, 0.0915601895333557, 
    0.00616280245499885, 0.0532923203114485, 0.0844405498056429, 
    0.0814661114083697, 0.00758389037765866, 0.0505124162741639, 
    0.0793622260623873, 0.0942666608574536, 0.108310199135366, 
    0.109488634410191, 0.0898656602609498, 0.0907137057391074, 
    0.128237505263251, 0.103704149471074, -0.0110309194845255, 
    0.259732769110997, 0.250043364839265, 0.0794164432441116, 
    -0.0478738498496144, 0.0588055274362479, 0.620842309888488, 
    0.264866098022939, -0.0829978637643982, 0.214378961238592, 
    0.541328581534837, 0.197300765319945, 0.0252196188537473, 
    -0.361527038264464, 0.683710125453051, 0.536091417178597, 
    -0.103988307152231, -0.507815284923747, 0.311630021193612, 
    0.359267754917219, -0.531831096465037, -0.130556595093433, 
    -0.155749810567491, -0.165466116535414, -0.209255780998915, 
    -0.123300878131894, -0.196956824129596, -0.150613684235885, 
    -0.191175071752558, -0.144271650657827, -0.19121196811559, 
    0.00355157055037347, -0.00446007885376627, 0.0452044391657172, 
    -0.00574042152878794, 0.0842167883088109, -0.00521847190544524, 
    0.0532425898127394, 0.0735126501108162, 0.093262878589597, 
    -0.0291241724067891, 0.0159914609085367, 0.148207487751391, 
    0.189090333095119, 0.139946650618642, 0.0972389314350417, 
    0.0928841522363968, 0.246099837435026, 0.32757324036514, 
    0.172393848153659, 0.0504702371772007, 0.434934301706619, 
    0.311331783053601, 0.0412138467775514, -0.0544519317886839, 
    0.675693723859732, 0.232111698550562, 0.027704433150273, 
    -0.100796926340485, 0.555372494424698, 0.290235804420846, 
    -0.0217675762936389, 0.414495701987367, 0.486218365720932, 
    0.14753043642684, 0.0125843358506638, -0.0769042567772465, 
    -0.342315510009786, 0.361448265617749, 0.387416355143108, 
    0.361520754248832, 0.447047747207461, 0.19952011896922, 
    0.0446477723677332, -0.0623931473612318, 0.137922766803976, 
    0.335186029417745, -0.180097893684538, -0.173615037722505, 
    -0.0650927611233991, 0.236812928345252, -0.0990258988617245, 
    -0.0560866487108668, -0.136885047621148, 0.00570237543912237, 
    -0.19936099574561, -0.00231735989688908, -0.424950851326741, 
    -0.120188194288667, -0.096669676691245, -0.328446582828074, 
    0.0071713250851265, 0.0999551182384014, 0.0639710642334791, 
    0.0797818664721054, 0.275846333985051, 0.287273427025843, 
    0.176470575920293, 0.135648754082377, 0.14345373298543, 
    0.220962700442482, 0.390303161687819, 0.274555003835145, 
    0.119243470569462, 0.403831516327363, 0.56173784066646, 
    0.227708839752995, -0.0306919263730219, 0.0884693999584852, 
    0.680762319915054, 0.274531270930891, 0.0713132339824379, 
    -0.0926398889648764, 0.722200604495818, 0.232092870884137, 
    -0.106992460733122, 0.220999170950093, 0.622273233034137, 
    0.0386635621812352, -0.613439325778759, 0.14190169801287, 
    0.720624214040383, 0.0198431513207834, -0.00183545845144248, 
    -0.0671039211515711, 0.448861976285388, 0.0732215641382952, 
    -0.440498616292869, 0.0899684176738192, 0.791044595922544, 
    0.450882124017497, 0.207610263706702, 0.240495797660992, 
    0.271450317700345, 0.270418978284899, 0.188381581188284, 
    0.0590261585833481, 0.146619951359807, 0.296858153234458, 
    -0.0411403822155674, 0.00560286312711974, -0.180851010941184, 
    0.558978521973957, 0.102179917634261, -0.181434143939867, 
    0.0395929880447385, 0.620299910132978, 0.0832046277536487, 
    0.0375317555098096, -0.221756702896113, -0.0459708614997093, 
    0.0479953103666063, 0.908427555076968, 0.292192093847985, 
    -0.265354879239894, 0.24219548005542, 0.612825985853963, 
    0.0820368645866223, 0.689989154086854, 0.590329688267019, 
    -0.0211461195923349, -0.0731846341894527, -0.243278329762208, 
    -0.055707083394738, -0.0560265005419407, -0.0915021574617694, 
    -0.0894224566577321, -0.0167187836453229, -0.129832807252423, 
    -0.00650878828568541, -0.114014481992152, 0.107787553931144, 
    0.16532613094685, 0.145534067673049, 0.14799552310357, 0.182790071414381, 
    0.112945425955457, 0.176654527225519, 0.365634102045627, 
    0.270065846628781, 0.116529679495494, 0.00962158044722199, 
    0.0464016922685072, -0.0196013904860974, 0.00634809369392168, 
    0.042171516040626, 0.00206275819189686, 0.0563632322719836, 
    0.0236765552626202, 0.0612910755050842, 0.0378333317296416, 
    0.0780991903089176, 0.0196404640822158, 0.0455790439404332, 
    0.0306610420173085, 0.035371378220429, 0.0347095001649931, 
    0.048880761618735, 0.0503351761107955, 0.0615969924131956, 
    0.00631046391961176, 0.0872779945370168, 0.104025995031339, 
    0.0941928364292851, 0.169715418739016, 0.204588347139586, 
    0.121164269918982, 0.112186433548382, 0.305863969627768, 
    0.17135646389182, -0.13392977522408, 0.210163718897646, 
    0.511614514985908, 0.1222624933486, -0.0119108579469744, 
    0.0679905345784401, -0.0533671900584977, 0.0738353822099579, 
    0.622650796247049, 0.524155238351818, 0.202459446959412, 
    0.0257052125645884, 0.620338770164126, 0.289022391856034, 
    0.119332833307705, 0.0747831474902381, 0.20037062201859, 
    -0.000266354122728268, 0.571412235538022, 0.336441062001593, 
    -0.0104763153115087,
  0.157502353400259, 0.145259237789725, 0.0310905882513193, 
    0.253536671038852, 0.224305991414814, 0.0107529224720935, 
    0.13367585492983, 0.301191346248993, 0.368224388470807, 
    0.407450029943979, -0.310630488727169, 0.614463801282197, 
    0.365716409487765, -0.35216973478414, 0.26659102140717, 
    0.735736975406582, -0.00231510661879163, -0.326329416336407, 
    1.04980877790163, 0.350317847801061, 0.115079726334113, 
    0.198039806400976, -0.0337606981703749, 0.137445029406771, 
    0.156353403346569, 0.197101193273172, 0.100741723657994, 
    -0.125148169454409, 0.153141759174166, 0.0508180615903279, 
    -0.221631610965388, 0.0526025865238598, -0.165896094946076, 
    0.0818776488829138, -0.317669394826484, -0.0455963219874539, 
    -0.205621952414434, -0.214459090722403, 0.11248186255878, 
    -0.242487657918407, 0.0535840637784843, 0.0121029600662749, 
    0.0374075823190001, 0.0318811304621744, 0.0543451246397773, 
    0.00220989381906739, 0.0195927832371665, 0.035035900116585, 
    0.0284330499675967, 0.000903564568417302, 0.000947082319184715, 
    0.219449334963012, 0.217728117784678, -0.017109586551245, 
    0.358392761210983, 0.370461552893536, 0.111611383876289, 
    0.0667037600813048, -0.00981962012948409, 0.244888169243617, 
    0.4535651166885, -0.390977000875098, 0.0529763230920226, 
    0.753780033379611, 0.321147652566676, 0.204264049841518, 
    0.636169998068147, 0.177274513865314, -0.495786207508714, 
    0.374400054659949, 0.671788983149915, 0.100068752380099, 
    -0.122060411733721, -0.200603235641632, -0.161354032951842, 
    -0.0824687454799961, -0.210969589119215, -0.125044311231615, 
    -0.139842978896043, -0.219151111641815, -0.0559829612795837, 
    -0.00764199627621055, -0.075132830154781, 0.000637386743425047, 
    -0.0827159227956754, -0.0212258477975538, -0.0569300321655585, 
    -0.048182492262415, 0.0417126684912341, -0.103940280250924, 
    0.0166052563345255, 0.0676984084794822, 0.0827399586856842, 
    0.059261926652809, 0.0634107910804208, 0.0685187454368488, 
    0.0654778545886736, 0.0789310046197017, 0.0669622300549718, 
    0.0290413911810329, 0.0790351231235987, 0.126693739698799, 
    0.171960550926792, 0.20711599064915, 0.176558378428779, 
    0.0720351609250164, 0.150361394909557, 0.439692825628241, 
    0.0679324920563681, -0.125339902493995, -0.136902235833898, 
    0.434089165161192, 0.352525501261006, 0.0820546118900363, 
    0.0402862608173843, 0.81197949667213, 0.286576757778727, 
    -0.0206234013801439, 0.220259890104761, 0.273598438866323, 
    -0.0576523851963089, 0.978441342302793, 0.490087407919691, 
    -0.0223999278914968, -0.204979023591916, 0.200294009190935, 
    0.267700475036603, 0.0294228685583529, 0.171046623304299, 
    0.0467302375160996, -0.424234252041651, -0.00762277459540701, 
    -0.21722608256542, -0.223489299716171, 0.0507827519831721, 
    -0.20930610735823, 0.070588419347148, -0.146056738767715, 
    0.00746272873863269, -0.207483540876034, -0.175238275525094, 
    0.192583430845057, 0.299026229126985, 0.039402022785265, 
    -0.0150302155983988, 0.663403987189962, 0.200188019421445, 
    -0.126801766961559, 0.0404321992853498, 0.581415408434701, 
    0.34069421228502, 0.178881113593016, 0.15857217361525, 0.204370237431509, 
    0.226403243415892, 0.176556446652212, 0.156562112102377, 
    0.204277033438779, 0.231244228579689, 0.180374009904231, 
    0.118099084763946, 0.10676887586318, 0.0985202121504863, 
    0.157021382101767, 0.180924535828524, 0.102690989007788, 
    0.114553940852504, 0.279638393007476, 0.161481670087747, 
    0.0748325270250039, 0.156736994604342, -0.116478200869401, 
    0.234103803219866, 0.623475758456424, 0.0124009293385995, 
    -0.0940000775701013, -0.148804149672211, 0.64912247023933, 
    0.112640015059164, -0.01618727261201, -0.16308952087993, 
    0.119563405030704, 0.614846518334007, 0.165020227752818, 
    0.034382982978914, -0.14992175288238, 0.546340380593565, 
    0.00139681032163795, -0.213495084757882, -0.1019588342095, 
    -0.220073690790921, -0.18532906103095, 0.0408374207566845, 
    -0.195280311483111, 0.0930479309542249, -0.0898273454326807, 
    0.116786257475138, -0.0795143350094983, 0.1400052138679, 
    -0.188229823716131, 0.108028972765991, 0.0749570204742467, 
    0.0788382645543679, 0.12093363699223, 0.130969416990369, 
    0.0917019139225718, 0.101741939600622, 0.130503619876512, 
    0.122516339551921, 0.0622668095992125, 0.095190034887865, 
    0.112404368511853, 0.142871813217396, 0.173630612293921, 
    0.128340908113812, 0.100975469632405, 0.262638255811351, 
    0.21841706381017, 0.0370863774899675, 0.0574480991363512, 
    -0.317657605717325, 0.292914648001159, 0.454317862880528, 
    0.0958042811103836, -0.0165498224135266, -0.234915115965905, 
    0.314647377451693, 0.448603751658645, 0.323447544036274, 
    0.179290760053694, -0.100325766674034, 0.000429321218165038, 
    0.299291043226289, 0.51422589514267, 0.208371320420568, 
    -0.104871784973436, 0.230006662515369, 0.309615187400173, 
    0.00777525842432786, -0.0737678689942043, -0.137165090588384, 
    -0.22550299248319, 0.0325420728907743, -0.089402697546319, 
    0.0575971941109137, -0.187641944702003, 0.0416039442787994, 
    -0.104216311420955, 0.0640170525956445, -0.250240075404957, 
    0.0187264188737506, 0.0867482825449755, 0.0670887784798834, 
    0.2641136660114, 0.263325629654317, 0.075451382197879, 0.232234340614766, 
    0.472091616766352, 0.197595575252325, -0.155869994791302, 
    0.755960565927498, 0.456836660641263, 0.146143689682296, 
    -0.367402495771815, 0.210399074745427, 0.811315669689133, 
    0.304662697469734, -0.18712713476887, 0.33810697439833, 0.52980378586849, 
    0.0916255832709449, 0.0403902295860892, -0.213462512777517, 
    0.00714587763099329, 0.406331845047809, 0.24080344755977, 
    0.111162386144701, 0.0199114410502799, 0.477925203663891, 
    0.100091120926845, -0.044740511802234, -0.0492385542802619, 
    -0.108053297988392, 0.0734581981936914, 0.103609243711531, 
    0.22704456659935, 0.222797078261167, -0.040918392782762, 
    -0.0358650571702389, -0.0257866571406131, 0.00402872787321369, 
    -0.155231909488706, 0.0528514064417575, -0.0296550553664035, 
    0.100377047643506, -0.109280802545725, 0.082308550175126, 
    -0.0494522979378258, 0.101055030466184, -0.191473012663139, 
    0.0498395054786607, 0.0569195950671343, 0.0685022715674447, 
    0.0615983087541711, 0.0643687265770248, 0.0612989307599404, 
    0.0698364442581749, 0.0976658839104068, 0.0876721252928047, 
    0.0048370640374424, 0.134645184896166, 0.179441969661397, 
    0.118323682694768, 0.0525065948482312, 0.105494550813954, 
    0.414931916216164, 0.220254139154481, -0.0409680949401552, 
    0.37837564283953, 0.241199181605709, -0.067478953246185, 
    0.0613147748423982, 0.466274615875983, 0.388980375217949, 
    0.202955125816898, 0.391583606570002, 0.769182562679005, 
    0.0432100703066311, -0.19903097108375, 0.197557760519723, 
    0.329406471824493, 0.00800822101832058, -0.0289156699924663, 
    0.0146262196427159, -0.051959196844613, 0.136779815008517, 
    0.11555315067342, -0.0647070964695453, -0.144220400006546, 
    0.220422890327365, -0.108440498215113, 0.226759872482911, 
    -0.202795766864345, 0.116293007580131, -0.167809453316842, 
    0.0963738150503614, -0.187842064424465, 0.0251412521456349, 
    -0.283334621875887, -0.12023976342078, -0.0208526355224582, 
    0.0424888393049131, 0.0132320329370938, 0.0253014911047841, 
    -0.0498436429047513, 0.00564502807235481, 0.00506045009450036, 
    0.0301630651977159, 0.0826029958451785, -0.0452728394122958,
  0.113110769374209, 0.243166229850663, 0.124045937323048, 0.054583301469879, 
    0.0301946554659302, -0.0650606142359442, 0.252063250630271, 
    0.169451982254627, 0.172526258609948, 0.118825683875398, 
    -0.0853829591963486, 0.0324852239502122, -0.00937221294176831, 
    0.0359261056413568, -0.27117379814703, -0.0161591275199414, 
    -0.181233663864512, -0.209979764317181, 0.166631179541857, 
    -0.251046680928404, -0.00293073649901894, 0.0672655637883789, 
    0.0775760518216286, 0.116800368580728, 0.14565035329223, 
    0.101411483903039, 0.0777796509935744, 0.158230207075626, 
    0.124861955533309, -0.00419449590095837, 0.123680351031997, 
    0.270656588973506, 0.229749677702297, 0.264867218399056, 
    0.257603719018213, 0.115297854673425, 0.267465829404279, 
    0.334339478642024, 0.254416589448641, 0.483766464089699, 
    0.547202204245315, 0.135729629414424, -0.418968520535672, 
    0.0628512004278401, 0.581663021738698, 0.21116209073552, 
    -0.2098778838739, 0.336486877788272, 0.475695578808955, 
    -0.138271658546793, -0.112812903357946, -0.192952575234122, 
    0.00458594890574515, -0.209984089037758, 0.0145867628588518, 
    -0.184441814139612, 0.0430852256923261, -0.157313411459811, 
    0.0648118885473285, -0.131452102453897, 0.122678302385078, 
    0.0528914221301492, 0.0756041462746023, 0.0785561003225847, 
    0.0940954025742263, 0.0724760157594302, 0.0960055437972073, 
    0.0703832399329389, 0.0812815110788469, 0.0384182772051752, 
    0.0467832806354465, 0.144950706192566, 0.130941115638466, 
    0.0744770192315197, 0.312372839779132, 0.233898075059678, 
    -0.00641715757119997, 0.449229820271319, 0.119529790961848, 
    -0.177097892448288, -0.193168931644284, -0.0554460731376378, 
    0.90463771914281, 0.405503639077015, -0.219220581032026, 
    0.268124055223572, 0.792950084106237, 0.325746465622542, 
    0.0860892979930153, 0.298143270912174, 0.267191370745152, 
    0.305441865614873, 0.210845467461338, 0.0593382704134989, 
    0.0121825763981069, -0.00602734293418722, 0.044610048696288, 
    0.0875757740009454, -0.0466870889137428, 0.0355766743446839, 
    0.0130475232446702, 0.0261297658170673, -0.37340494561719, 
    -0.0368024489266082, -0.101045076432251, -0.258239929767087, 
    0.0793788095780935, -0.0510666909739416, 0.0907095282831738, 
    -0.215651144963645, 0.0206473216259914, 0.00665509402916334, 
    0.0149978615098757, 0.0100986033830034, 0.0145974733965707, 
    0.00621760062819776, -0.0391799011037446, 0.107650763846851, 
    0.232640843098582, -0.248323660714152, 0.359910205857907, 
    0.308283130648033, -0.0403016296800818, 0.266094136358412, 
    0.443800483396529, 0.102909269407645, 0.00205505347979712, 
    0.518196360317461, 0.560601065148747, 0.362970061189523, 
    -0.172841529114916, 0.476374856013119, 0.19368876141308, 
    0.653873646185944, 0.916112654542603, -0.197627643837376, 
    -0.537897677764344, 0.450225049864194, -0.0600866347263088, 
    -0.432150566925117, -0.304360333783805, -0.0479716393583148, 
    -0.268646855655731, -0.227086376926581, 0.0700623168231607, 
    -0.263293257756073, 0.119317578323161, -0.197437213075384, 
    0.076178774154549, -0.253108215105615, 0.0422737601654088, 
    0.12054108059113, 0.136641750680392, 0.210421044949623, 
    0.186783629593375, 0.13905753746566, 0.144848112554478, 
    0.192327695836824, 0.168076475554735, 0.149374640050117, 
    0.170210386529552, 0.183805466916627, 0.171927472321783, 
    0.176894203650901, 0.194864280690174, 0.173530679489964, 
    0.130768865406163, 0.139729014276302, 0.20480933247203, 
    0.201977865164631, 0.132936345190578, 0.112985567649379, 
    0.111903608167299, 0.114548005019457, 0.122983634573303, 
    0.106423388365733, 0.110583014699078, 0.151583500019278, 
    0.126226411163027, 0.0553600922703435, 0.154595183911299, 
    0.238037289988047, 0.154990961059473, 0.0518016944022323, 
    0.263749110561088, 0.381594301726216, 0.161764188866372, 
    -0.0531759385032835, 0.126193528675732, 0.584949948842059, 
    0.129227189602888, -0.166141128916104, 0.0279592398417646, 
    0.548214711874066, 0.19231900921639, 0.161133771721255, 
    -0.136820775093561, 0.451209055312952, 0.304674817514515, 
    0.167780517190589, 0.295521574652793, 0.270876158353172, 
    -0.22474533360098, 0.0738500130786763, 0.579806786967743, 
    0.534660232709005, 0.108978451526543, -0.193030982440631, 
    -0.0307483414827377, 0.0272075751216836, 0.393996608078313, 
    0.443506111392713, 0.0312565226626866, -0.0613266805849638, 
    -0.0317420567617301, 0.219610466075036, 0.15781854754785, 
    0.0441687996590385, -0.104408539397697, -0.109907682925413, 
    -0.277658134245441, 0.0327433303905064, -0.318563207174062, 
    -0.143936191174706, -0.162042030244665, -0.200061825423529, 
    -0.119636173042692, -0.182972403394752, -0.0437351962755151, 
    -0.182553251774956, -0.00058678961248114, 0.055977718039046, 
    0.0617031494891923, 0.0718104704136014, 0.0869361108540848, 
    0.0508570435892655, 0.0368705165419777, 0.117701487359818, 
    0.0748496722923496, 0.0482702297864364, 0.202754283975821, 
    -0.0739015492240094, 0.103456899826072, 0.284744452934465, 
    0.5534368207949, 0.356806007852205, 0.0530079199282562, 
    0.513184191350424, 0.350496601310196, 0.0463073283558085, 
    -0.443442869012365, -0.0484056049184182, 0.664219373492727, 
    0.158793648271918, 0.078039320646701, -0.449542864060294, 
    0.32266163005172, 0.6788791510365, -0.253451211606244, 
    0.00577190413784564, -0.330271046494349, 0.0180653036602235, 
    -0.161393897497847, -0.168036828915241, -0.0187540819109256, 
    -0.185948976253649, -0.00995135780889837, -0.153609689734421, 
    0.0166245229516392, -0.165466611007157, 0.0576709604574617, 
    0.0877925578019883, 0.12678327368176, 0.183896129357965, 
    0.26383856163845, 0.316184131923753, 0.235707488398262, 
    0.130097822413376, 0.219207923128678, 0.369816963559706, 
    0.295941993588743, 0.204537422152366, 0.173555084695168, 
    0.190103414627083, 0.202805635478494, 0.172541133101736, 
    0.153950499374714, 0.190362138524883, 0.213675755094604, 
    0.193129289038727, 0.144076280286127, 0.0687970602198445, 
    0.281316962686943, 0.324160947848992, 0.116165232404399, 
    -0.0697429991647865, 0.30837003432648, 0.462221576314684, 
    0.127330268420469, -0.188287505039642, 0.0109931886721591, 
    0.360663973907642, 0.509482491954241, 0.282400589574362, 
    -0.205287848028388, 0.40578643379195, 0.302181979706903, 
    -0.0394788244895361, 0.217240228576676, 0.51599568369717, 
    0.0499459192637028, -0.0136394207497576, 0.140301076335918, 
    0.108648231280715, -0.110295761600352, 0.125661237161031, 
    0.142262943403419, 0.0269692864010681, 0.00313165039403407, 
    -0.022386694630649, 0.0516477861130861, -0.246787785871744, 
    0.0883829528711807, -0.23682104037986, -0.077974009831981, 
    -0.106939959151434, -0.0102419120854577, -0.0904571038072826, 
    0.0294805638075325, -0.275429140060868, -0.0523859489683905, 
    0.0763600582707453, 0.0944855805791494, 0.0611935504141765, 
    0.133746711889194, 0.191509047091194, 0.158139491687947, 
    0.178833812680344, 0.208570112951671, 0.160431202577556, 
    0.135054327417448, -0.0466311369685508, 0.453443376642802, 
    0.490696195838725, 0.14909253000501, -0.221712585572185, 
    0.33000510651747, 0.565220490266394, 0.0811110570327767, 
    -0.131540769244073, -0.0884351615452937, 0.437763262513218, 
    0.350329776291159, 0.218666680263082, 0.247066379044243, 
    0.200878119668319, -0.344846551574494, 0.325324843305502, 
    0.490692560512325, 0.205705515533692,
  -0.0171799611553433, -0.149149831214316, 0.0526067298803594, 
    -0.062901988190245, 0.0379189806845856, -0.140048246295343, 
    0.011941449527631, -0.0639175837486518, -0.00683517101832853, 
    -0.154326233631211, -0.0595884271428034, 0.0227563990741852, 
    0.207719369165313, 0.238839192656601, 0.0738416495779681, 
    -0.168073523217583, 0.0332967682136856, 0.391857149918082, 
    0.198390246925333, 0.374062538471783, -0.29113248329807, 
    0.402669826717691, 0.47396560064846, 0.467629198551566, 
    0.286236343131944, -0.175049904378945, 0.184296696469614, 
    0.288911169906486, 0.148891718075379, 0.841964187604242, 
    0.64165328247309, 0.219531005963, 0.0798573606855314, 
    -0.0233552749976337, 0.190081109357216, 0.361408689236928, 
    -0.133799000575022, -0.134202000721263, 0.135272149861692, 
    0.186698659594406, -0.253174344322953, -0.106764151995352, 
    -0.13757307506734, -0.142622598718481, -0.10111939650371, 
    -0.158057642314779, -0.0867527395896094, -0.223059202049689, 
    -0.0509689148344903, -0.137559329027693, -0.0652264802152339, 
    0.025741853775242, 0.0490782665991174, 0.0594219618919824, 
    -0.088184782035781, 0.0572218037845262, -0.0779593597594693, 
    -0.0141934185480121, -0.0278663422165143, 0.0125535860997625, 
    -0.0397474183419094, 0.0270378794006251, 0.146818197013589, 
    0.101613729971159, 0.229906602940589, 0.225156766474334, 
    0.0169453336414703, 0.0463734925111536, 0.545473687101933, 
    0.249814750870603, -0.157526532995344, -0.0554126617937781, 
    0.893555293335575, 0.517963041282439, 0.0310563158613352, 
    -0.184178430451259, 0.0852727773865347, -0.741642933656504, 
    -0.163029409295066, 0.786536023800582, -0.24198790198095, 
    -0.17362060577695, -0.181515451458828, -0.0732546262260028, 
    -0.171867662878737, -0.1173972182267, -0.00010168337283549, 
    -0.142473437122681, 0.0421936517650969, -0.114858946826361, 
    0.0599460930456831, 0.067866133421753, 0.124592373061543, 
    -0.00758156561087385, 0.0547824124634355, 0.0206634713365632, 
    0.0301898878573724, 0.0508901339558479, 0.0646466213441116, 
    0.135886112007218, -0.0145596189204573, 0.0550459241116978, 
    0.0002861202875101, 0.0142795589064162, -0.0709552743958867, 
    -0.00348466590915066, 0.00666082510031461, 0.0114691041151246, 
    0.0651219928374858, -0.0390764412445087, 0.030962716324424, 
    0.0455343334013282, 0.0466296048570963, 0.0465846319553452, 
    0.052442459716531, 0.0583466278271453, 0.0412041811373394, 
    0.0105406860864324, 0.059425070807307, 0.156121618855109, 
    -0.263012029792867, 0.595696617511244, 0.406724487232802, 
    -0.237362590344905, 0.188988979689067, 0.777985861711284, 
    0.198463340064151, 0.15548069849582, 0.00612942054631557, 
    -0.423295123166903, 0.648864331975652, 0.642176335279691, 
    0.287028133371644, -0.104433704150175, 0.136723985480888, 
    -0.0069939571499687, 1.20556949938343, 0.399099293364301, 
    -0.0279714340463824, 0.724155686174536, 0.385277661609954, 
    0.00776346144046851, -0.0467036425475285, -0.0491033883032346, 
    -0.108356906407949, 0.117663218486584, 0.00499062155848493, 
    -0.155858668797763, 0.063129822987931, 0.0828940465063095, 
    -0.0126527858935498, -0.0903832023991425, 0.462088486490115, 
    0.253375484204782, 0.115535168410348, -0.177896733510283, 
    0.103168643855702, 0.402221002476501, 0.0857925840804605, 
    0.0421140403209127, 0.0842887753124396, -0.0512291484322296, 
    0.579850581503569, 0.0716509012601754, -0.0155284393395433, 
    -0.103252724204972, 0.505843451778101, 0.191576274598644, 
    -0.0885767908896117, 0.509054285601304, 0.43872594270355, 
    0.205359720163107, 0.134631560396753, 0.125202292469402, 
    0.121735441794083, 0.116866054089072, 0.156320519405999, 
    0.141221136075708, 0.00315472355713423, 0.0679210510154102, 
    0.346649641457932, 0.305751260480562, 0.238618787338389, 
    -0.155997524591776, 0.378617408241208, 0.294858259812392, 
    0.0532754228556452, 0.381515833380599, 0.35806327265903, 
    -0.0292216055068466, 0.0143273539354631, 0.632385060038127, 
    0.204083251850681, -0.0998164180506859, 0.397189859986729, 
    0.418573355126848, 0.132548811617371, 0.0612198976296153, 
    0.530580620425079, 0.177075858182651, -0.0156566181786078, 
    0.00899745406710961, -0.0301042787177528, -0.012445550998315, 
    0.00629494768596625, -0.0182759088004021, 0.00532327476455991, 
    0.00700145596878393, 0.0320557385806308, 0.0688284019448204, 
    -0.121421415410833, 0.254369448896725, 0.260435607143342, 
    0.0615423660655272, 0.0222013851973474, -0.0559649724436832, 
    0.296261693093028, 0.492735305239845, 0.231875172505135, 
    0.166806766623921, 0.0655212727174421, 0.767246099229508, 
    0.0808732253133787, 0.0771458266105206, -0.274428581577782, 
    0.114314851261003, 0.682063258425041, 0.406249699130616, 
    0.0248839061190097, 0.576447146056333, 0.273013910490554, 
    0.0505861450279557, 0.21051207547556, 0.321318459004436, 
    0.23727840968426, 0.117085605224456, -0.150216209056891, 
    0.285301069595528, 0.105244154939212, -0.213827270515877, 
    -0.0184867467045809, -0.203998759955438, -0.00130156822829261, 
    -0.245478368916458, -0.127134178096418, -0.0979147206513284, 
    -0.12207144532645, 0.0348123827435666, -0.123103181143431, 
    0.0246479032282438, -0.0519171914724182, 0.0755771046139758, 
    -0.0195019744736955, 0.0678871647673321, -0.0134022398489127, 
    0.058955332940524, -0.105389088098278, 0.00429297784619848, 
    -0.0595503091802933, -0.066357823201383, 0.0222992456725434, 
    0.0529159115538329, 0.0875855975386287, 0.0915454574462845, 
    0.0802272250581911, 0.0793650158877437, 0.0731324163435948, 
    0.112023028981017, 0.102264008096496, -0.0612679619131553, 
    0.285944182452857, 0.263902031766028, 0.0302240540554396, 
    0.134822875137616, 0.188029215570959, 0.271790694211657, 
    0.584908598685445, 0.410279706450668, 0.165606565062829, 
    0.0695420814321664, -0.0786215030914595, 0.0494983823387708, 
    -0.346715127715628, 0.695333398108679, 0.449532606362227, 
    0.301807322678377, 0.666490673492928, 0.178736743100003, 
    0.0932820287073474, 0.172888369444521, -0.347308914114575, 
    -0.205856349521554, 0.0537341531493522, -0.142444703470103, 
    0.157071245364844, -0.189205207479311, 0.127189168242341, 
    -0.237321116647459, 0.0601580824638877, -0.223887586215347, 
    0.010004390951283, 0.0944921027738885, 0.135953300692838, 
    0.173747476470793, 0.209424656667874, 0.228040424373826, 
    0.23260992811397, 0.233419739974765, 0.201606855403617, 
    0.175800109436945, 0.157809368424511, 0.170234742040323, 
    0.176849764077255, 0.180330576235746, 0.184720167961402, 
    0.166479092305044, 0.165176647902241, 0.206624075998241, 
    0.208248630815811, 0.173076272916259, 0.167752815773998, 
    0.175387978611574, 0.181705313736955, 0.206954217945695, 
    0.191234680288564, 0.160782631088823, 0.290264698224961, 
    0.333204060928206, 0.149230901068534, -0.016399965638866, 
    0.523870179213817, 0.259371276841683, -0.0131562682527517, 
    0.0248044156968364, 0.551437724448263, 0.232592622972349, 
    0.119454114697646, -0.202999803583719, 0.117418436395951, 
    0.402655841424923, 0.419538949080774, 0.195710390371801, 
    -0.147833623294695, 0.202367748818159, 0.132731059234796, 
    0.20375135149467, 0.778124784964752, 0.309671111365116, 
    0.0543757479930625, 0.257551250959572, 0.272940138304141, 
    -0.0804695311401996, -0.146796854145558, 0.0721299712215468, 
    0.114441252701485, -0.0345506977657104, 0.14824717131163, 
    0.122261104124739, -0.0347780946374042, -0.0543812074793684,
  0.0515586930619908, -0.101576046891299, 0.0193458695226999, 
    -0.00548025752506112, 0.0283135543271324, -0.119085332412687, 
    0.0161959224989158, -0.03535090926484, 0.00921411470960523, 
    -0.0951395562928867, 0.018349993176248, -0.0277783660492999, 
    0.061966979620343, 0.125268573742425, 0.0533846169761896, 
    0.0015560647156528, 0.0487480296162853, 0.218050809663101, 
    -0.128953108903098, -0.264055691468015, -0.110251912084424, 
    0.685555976399041, -0.687671454658813, -0.545417909959208, 
    -0.540973723902162, 0.383937957763206, 0.847121841418448, 
    0.489055545439348, -0.0879383265672431, 0.981240943518228, 
    0.415176222290105, 0.113922430673121, 0.176430694085219, 
    0.336809700996446, 0.121127951089054, 0.28246746084069, 
    0.266028832823219, 0.0493243353246152, 0.341710841864261, 
    0.228019853765242, -0.166121362648993, -0.0809311434988559, 
    -0.133896605334635, -0.0807894604025116, -0.193680981736912, 
    -0.116571694028008, -0.0125064938522723, -0.0866776589937674, 
    0.0772248876808906, -0.236117952631221, 0.101620600964505, 
    0.186114192296016, 0.0486598748936772, -0.0342553499719982, 
    -0.045281523790776, 0.433120465685626, 0.450480683471756, 
    0.11385433828592, -0.0896321371809352, 0.0364293532372991, 
    0.294389189478563, 0.27294297690625, 0.190962644843421, 
    0.145225546505394, 0.142461937454165, 0.159486941782646, 
    0.15335060719223, 0.155475954215864, 0.16743695089402, 0.164219764032161, 
    0.132374651626847, 0.109071068893089, 0.0979569302316973, 
    0.110118679678369, 0.1740831392126, 0.223767592045861, 0.185129691300088, 
    0.129118406554732, 0.122188219975067, 0.160635553476194, 
    0.204539944841522, 0.214746608554602, 0.201541024283611, 
    0.184759173212996, 0.165789333532498, 0.140365456886035, 
    0.152313677833162, 0.19803325755997, 0.166313014323525, 
    0.141974088100663, 0.267885445219774, 0.218069698322822, 
    0.0520780007993309, 0.121026469827469, 0.454525154563453, 
    0.243494432840287, 0.0567499856963541, -0.0698583128344704, 
    0.274445040966174, 0.408993864199777, 0.285835179783819, 
    0.0948940893910154, -0.18799096082774, -0.0231052436106799, 
    0.383548829534688, 0.496809507188931, 0.322358248957014, 
    -0.00661231252903724, 0.512064182690934, 0.68621626340151, 
    -0.249374063561183, -0.246908436747863, 0.00680215502634238, 
    0.4424755134183, 0.0077442206473439, -0.278818146988527, 
    0.33715875001119, 0.381925372413133, -0.20326951230283, 
    -0.0266880600240196, -0.508785464782717, -0.177758897807782, 
    -0.280779018098283, -0.290585994232657, -0.195709682089403, 
    -0.248705057062569, -0.0295266252601117, -0.215644136291406, 
    0.214085876250975, -0.261399493667067, 0.159570686604642, 
    0.0363350385592889, 0.0642831226895387, 0.0792414309408872, 
    0.0796965151247939, 0.0266265870734565, 0.020381420612009, 
    0.0997053314576563, 0.102423175459203, 0.0195128601954312, 
    0.084781270379774, 0.107466277627943, 0.106000372163496, 
    0.130075787894118, 0.0776166857136681, 0.0874499561084303, 
    0.245684535535704, 0.0727622453126801, 0.121404965103154, 
    -0.101036588552284, 0.817671591451781, -0.173345158104585, 
    -0.492189149779992, -0.101191793385409, 0.718239035560708, 
    0.434997155976577, 0.208621538371328, 0.0967924536942338, 
    0.017035618481705, -0.30686546532265, -0.0429603086219748, 
    0.46661950424968, 0.281930424230819, 0.150680808268877, 
    0.151312947499337, 0.151358792373709, 0.112633774791049, 
    0.100420608403123, 0.125730104299242, 0.130297298378911, 
    0.119145211017802, 0.112492561812731, 0.103196836756781, 
    0.119186671054732, 0.146950303874655, 0.115129015399984, 
    0.0714338916151676, 0.0826678058042333, 0.0505565679214854, 
    0.237402046316764, 0.319738839594594, 0.0478905588356109, 
    -0.125100373594233, 0.0892665011948989, 0.747845026096695, 
    0.01640357453822, -0.0191441070423385, -0.276308672986621, 
    0.340526648057914, 0.486264228206763, 0.0161895658026918, 
    -0.259139411081462, -0.101757392335887, 0.488541855005929, 
    0.0986704168478521, 0.0392222316162908, 0.0456320375848321, 
    0.0230730660653914, 0.609414911123059, -0.0238869701016543, 
    -0.150300509892579, -0.0110247470111617, -0.115361881397087, 
    0.0108290781775326, 0.00750124670765473, 0.118766163199887, 
    -0.135770385136095, 0.0213338917315314, 0.0863088055347944, 
    -0.166494758671056, 0.461799275676106, 0.0959677761308932, 
    -0.0515278934122586, 0.467102069972723, 0.410304730599963, 
    0.21310670962515, 0.184817829151324, 0.14517607869801, 
    -0.0889752881484587, -0.201502700941096, 0.861926736129978, 
    -0.0289921054560541, -0.46213584259934, 0.0555245287733048, 
    0.700558558812917, 0.302657821306245, 0.39454631867605, 
    -0.0570390726381627, 0.721915295588121, 0.249742759482605, 
    -0.0138876849803416, -0.312048074193977, -0.0126909570860555, 
    0.394718987272217, 0.123408886716012, 0.086007485978007, 
    -0.164269369305667, 0.306974727202738, 0.193728926683596, 
    -0.0602090752616265, 0.304882154947019, 0.28065415224519, 
    0.0423862777960092, -0.17322722369907, 0.336413782708595, 
    0.359736360864696, 0.119333625632006, 0.0160753784806321, 
    -0.0803717447880907, -0.173971369679842, 0.295918910794819, 
    0.329297963378183, 0.136995812430984, -0.110082677034769, 
    0.211789761121343, 0.367006141737399, 0.11363925191991, 
    -0.0214549250839233, -0.082807974384196, 0.343438089183498, 
    0.392898699004098, 0.384936729868372, 0.254718308294157, 
    -0.196329044551938, 0.28948422229302, 0.378422656886208, 
    0.0856566162061873, 0.256297787146701, 0.476500909855989, 
    0.239841490337767, 0.273374773273147, 0.365241424796392, 
    -0.113520363167592, 0.298407763595393, 0.709005056164838, 
    0.0246704968198962, -0.128849513402225, 0.160298949836923, 
    0.365760111592875, -0.00673628061161408, -0.0958401359156908, 
    0.0337027321868472, -0.0751898358993612, 0.0219869439551741, 
    -0.124686067453978, -0.025555035440284, -0.0508114172007494, 
    -0.0507312344134224, 0.12546264116755, -0.14631763881743, 
    0.10765515085646, 0.213368772896783, 0.0259791358533799, 
    0.271406127913053, 0.229265247168354, 0.237746437563642, 
    0.503791904033291, 0.140852358363188, -0.00687451061801764, 
    -0.242099453304264, 0.123114101058278, 0.553389564053252, 
    -0.00218764811156766, 0.557000262952399, 0.877656143113579, 
    0.524642384764004, 0.110706310629109, -0.222331484469281, 
    -0.173084965245345, 0.128826100056706, 0.57851618735544, 
    0.286103249044374, -0.0813658706134464, -0.032161170652289, 
    -0.0946460605857763, 0.245318995538973, -0.0924017864643038, 
    0.0553025258163135, 0.102885841207767, -0.0817450597824521, 
    0.169282991460704, -0.22412096062789, 0.187340082892526, 
    -0.202515744067264, 0.134933997881211, -0.165118853424037, 
    0.12979593550768, -0.14968064200219, 0.0857862004888571, 
    -0.263511397266487, -0.0408039120663773, 0.0487186117268787, 
    0.03807965037783, 0.122810854680574, 0.0866262742544439, 
    0.0847277496160915, 0.297356276165316, 0.0859514847261473, 
    -0.0322840836149602, 0.0102410068572889, 0.662473337175815, 
    0.0322244930891414, 0.0545292903629348, -0.19465590912654, 
    -0.206836954365366, 0.90212199995021, -0.0526279322219945, 
    -0.27423612786842, 0.296996115732209, 0.35092744528162, 
    -0.210206055054661, -0.103749146410652, -0.00368566302593128, 
    0.0065251263533774, -0.0748374937368756, -0.0611586922666073, 
    -0.0466249338673776, -0.0381454526555834, -0.0895148408647864, 
    -0.0817910322242549,
  0.227411156628522, 0.724476495571169, 0.303812372322544, 
    0.0569471314258069, -0.295230997197926, 0.0578245702039361, 
    0.540336180971636, 0.330054354363666, 0.181020925261158, 
    0.106488490637398, -0.0759380815534723, -0.0191483087935618, 
    -0.0692086248686177, 0.171720437422543, 0.0136859322404053, 
    -0.0891578029754158, 0.0360258483478808, -0.00172290374511178, 
    -0.172527827156402, -0.094381026839027, -0.0273444429396408, 
    -0.00563587021164715, 0.0211136377569534, -0.00941852326362361, 
    0.0512858276701189, -0.00584173293458694, -0.0412966192922729, 
    0.118024934558021, 0.0848030478714258, -0.0647783742578345, 
    -0.221910892753625, 0.0676036266027085, 0.437303994319183, 
    0.347263664728918, 0.182965027364632, -0.180395492110958, 
    0.241554540919126, 0.427308236837243, 0.357848318651801, 
    0.0896383152729396, -0.275255089366694, -0.0691839917974987, 
    0.632860280101617, 0.180290434113507, 0.0239029489739134, 
    -0.0565561005844757, 0.23586623394531, 1.0977046954058, 0.80467187541932, 
    0.228182961609973, -0.0882548243474644, 0.42410890862758, 
    0.357300943224534, 0.0496423693021987, -0.0662679280715083, 
    0.163123612546188, 0.0547775352587948, -0.025387563386452, 
    -0.0207788029760014, -0.0543501771483188, -0.00104108180477566, 
    -0.105632456232276, 0.0165103626171048, 0.132018292800827, 
    -0.0106831920661713, -0.0740163419538472, 0.0286566693031883, 
    -0.114166493094355, 0.0827982557967728, -0.0672924755557082, 
    -0.127528265812346, -0.0517392229341372, -0.051498467340099, 
    -0.0199747416141795, -0.0403829645261592, 0.0496108987120049, 
    -0.296794598587657, 0.0300706481756901, -0.17152475325456, 
    -0.139689467606323, -0.0104218560172127, 0.0269753891271798, 
    0.09295242304578, 0.123311772563098, 0.109199383938144, 
    0.0856107934148412, 0.0714764562728191, 0.130206900628702, 
    0.111630701642098, 0.00818545540587214, 0.109539896578165, 
    0.314502151407176, 0.235975961285068, 0.0606197496318931, 
    0.0553587065797627, 0.457859327873036, 0.393531046845342, 
    0.130703309966039, -0.231776228638036, 0.23659500068647, 
    0.541583256733991, 0.0832172565101358, -0.055560820438714, 
    -0.196180213279414, 0.416884591821492, 0.474215118349344, 
    0.207838562115592, -0.153989638550276, 0.304136397774358, 
    0.400952988590536, 0.290982790911194, 0.238833415832372, 
    -0.0358474667254793, 0.495267847671719, 0.180712233206882, 
    0.0442828920167183, 0.127174018991244, -0.048066631535687, 
    0.107221085456183, 0.706216739951781, 0.086811736243572, 
    -0.0511403086027902, -0.04003532536142, -0.00882928174347823, 
    -0.0651752917492541, -0.00813415979994451, -0.0578457887502119, 
    -0.193607476831391, -0.102553483435725, -0.13585878882572, 
    -0.124164584605176, -0.143218553777946, -0.0197393811949466, 
    -0.154324136134934, 0.0276335064876238, -0.130883209882545, 
    0.0461735049423616, -0.057327182815143, 0.0913007295460941, 
    -0.131481368805984, 0.033001733311741, 0.0596899398282287, 
    0.0691197747239519, 0.0711477627326754, 0.0751717242738202, 
    0.0609449914742296, 0.0619421074978749, 0.102320149435308, 
    0.0890136361009418, -0.0323532316179334, 0.184174650620676, 
    0.229026869317043, 0.0918776950213912, 0.138498586343853, 
    0.346030436877073, 0.22343963444424, 0.0953567098495499, 
    0.302756510569354, 0.302038385720401, 0.0124641412725657, 
    0.164428232595675, 0.684221443692899, 0.255889109456796, 
    0.119151653868524, 0.385694910528948, -0.0737018372733952, 
    -0.064149783740448, -0.513465475409255, 0.0482391460254489, 
    0.421860169426446, -0.255427930181711, 0.0631996657878874, 
    -0.198450212652675, -0.0405825809860714, -0.186868169183442, 
    -0.052093599050898, -0.190746580968184, -0.114519988233562, 
    -0.0741439575989148, -0.197393945683697, 0.0653058426286391, 
    0.0350840418666565, 0.00468420898963108, 0.00886231118761979, 
    -0.012311050403055, -0.0602300007398513, 0.0489842567690429, 
    0.0769055707005749, 0.0737930331724731, -0.0206961405202172, 
    0.0288644939424314, 0.0787877261213989, 0.107707413161196, 
    0.135339604447053, 0.151995642710653, 0.121615362118167, 
    0.112935128287359, 0.183002845016636, 0.172731875034107, 
    0.113799522614905, 0.11179733058747, 0.0387210691516236, 
    0.320132630194124, 0.432787296763491, 0.141671080799713, 
    -0.161135373668136, 0.122978193286887, 0.610137685533648, 
    0.142422311547361, -0.149524521805098, 0.262422770235782, 
    0.317637096505481, -0.0135646093520388, 0.568723486766334, 
    0.587664122261861, 0.0627671591967922, -0.251432563711999, 
    0.101470838156494, 0.499631196482187, 0.168822617002731, 
    0.0376835372793113, -0.180733094775059, 0.24220273834028, 
    0.0652028609300039, -0.0606227132113185, 0.0940053071562737, 
    0.201466394019784, -0.111810023911469, -0.0966706786242274, 
    -0.0109736901819546, -0.334724522115788, -0.210509472637818, 
    0.0911252694911503, -0.120799762054803, 0.166950469325691, 
    -0.179149391752723, 0.00943704786697398, -0.0565250156183373, 
    0.077120981929537, -0.221144389054981, 0.0548432942803197, 
    0.0639333902134932, 0.070008757995584, 0.0496515972840183, 
    0.0576847916401782, 0.0200684064584239, 0.0467758201501477, 
    0.0367647980052136, 0.031417068506687, 0.0321363824856502, 
    0.0961308817086435, 0.0771959621529841, 0.110074289557941, 
    0.180300125254476, 0.206082407660932, 0.198607713537784, 
    0.196082548231344, 0.234872957409535, 0.180941932588854, 
    -0.317434895501519, 0.269040247075639, 0.356400261504367, 
    0.0313218441610145, 0.660843729362756, 0.613931029430702, 
    0.251498275214197, 0.174167994517862, 0.238676458710445, 
    -0.0546253118829521, 0.418431952912979, 0.572812448303319, 
    0.123019186646898, -0.0293151990100152, -0.0779009756762058, 
    0.0701924780102495, -0.0499805548956437, -0.106111578710284, 
    0.000726909957729754, -0.0741921942970192, -0.0396387439121407, 
    0.0496883981036658, -0.168245686215908, 0.129615014339435, 
    -0.170619720784693, 0.00468566157887237, -0.188742926800034, 
    -0.0369456994025923, -0.105708264222555, -0.0198938393924779, 
    -0.229650326100938, -0.0559944516772143, 0.0473773481385661, 
    0.194816676610088, 0.179931931004587, 0.105887542027708, 
    0.113274932846837, 0.198723902497842, 0.270055252452657, 
    0.269865137683374, 0.198404242326467, 0.168505352954545, 
    0.182651812538081, 0.142912376280145, 0.162409164855611, 
    0.204168486889047, 0.199474228190234, 0.060703893138552, 
    -0.0704934262334823, 0.0972365176480152, 0.191618234637908, 
    0.272039388318037, 0.379520981480088, 0.181498122591008, 
    -0.137566094376819, 1.02802942826268, 0.406874068991443, 
    0.0960434876743859, 0.224214007201693, -0.32886821651415, 
    0.231703633147608, 0.332149935218027, 0.189490173694523, 
    0.0744871642138687, 0.0956943378680137, 0.281512554349861, 
    -0.0474661522492589, -0.113365172400051, 0.12099986402785, 
    0.0115915086259852, -0.0587230733933553, -0.238948307154524, 
    0.0615437885342805, -0.142155205114786, 0.0321361514537108, 
    -0.360516907211299, -0.0596660098926855, -0.125772855496705, 
    -0.22087639131189, 0.152659505674906, -0.29717623924312, 
    -0.0588163375210619, 0.0632510692490067, 0.0450923075613694, 
    0.113088513638308, 0.170173535546616, 0.0554859809461335, 
    0.0550620256417234, 0.235110104449056, 0.318675342992256, 
    0.309104691453773, -0.110935373876259, 0.646479189149153, 
    0.308281868318187, -0.0870125328038221, 0.446923074116469, 
    0.47532485355906, 0.101712098074, -0.360304344205196, 0.710747225118693, 
    0.399290186130916,
  0.00899532861534329, 0.0487698436989483, 0.174003152197788, 
    0.148109657472154, 0.0669178205199174, -0.0175380748215986, 
    0.155940187374345, 0.231199958684225, 0.234922206169297, 
    0.0755482531938434, -0.088000252800137, -0.194061650577173, 
    0.587017123838912, 0.207778657215605, 0.0708200882872045, 
    -0.223604316278056, 0.0294809960987856, 0.428632873364933, 
    0.355462970008355, 0.432973507286222, 0.324905019019537, 
    -0.00816284581807003, -0.0888609520978455, 0.0681271264536712, 
    -0.00372695711435103, 0.258128101345899, -0.0733602305440787, 
    -0.0418364197881616, 0.00884527264071122, -0.0112588258309983, 
    -0.0604874752237512, -0.174231337926308, -0.0405850866123951, 
    -0.0792225831107922, -0.0194520301050009, -0.273957612593407, 
    0.0108516876951311, -0.161511298504965, -0.0106791536311708, 
    -0.294387899351056, -0.0344768919818771, 0.0232167942886722, 
    0.120248645321409, 0.132293941330484, 0.108937405028993, 
    0.135015722092499, 0.176168903656721, 0.184245126109879, 
    0.143588563153016, 0.0925301090054042, 0.175796567858196, 
    0.195547514046721, 0.237765305406825, 0.383858088453301, 
    0.329158963309999, 0.132862789450928, 0.104112795553418, 
    0.483450337346063, 0.385928472384899, 0.238151725786832, 
    0.151277815513988, -0.178552294815203, -0.114433058349348, 
    0.491182560206956, 0.226190013327854, -0.172554201015886, 
    0.662712509241629, 0.762532237571008, 0.21269050735109, 
    0.00740592948667955, -0.0987737900090397, 0.280194007287511, 
    0.11231390463293, 0.019128526144106, 0.0342624873757158, 
    0.12745329670938, 0.0556868065556163, -0.0301465015726798, 
    0.123852170270206, 0.135701032519582, 0.0651417044203854, 
    0.0457975652615327, 0.0472496953092126, 0.0446213006335089, 
    0.0499373339671355, 0.0383326286672276, 0.0230809507408953, 
    0.102757231703493, 0.0391066649577344, -0.0182569356816303, 
    -0.149575073266776, 0.268369386261483, 0.441821474733111, 
    0.258452061145332, -0.259040290581012, 0.334548620186376, 
    0.457064376671845, 0.148284582245683, 0.0160321548763003, 
    0.0136583355924093, 0.272756446716933, 0.054234570990058, 
    0.963893119027579, 0.508181357023742, -0.0389776173990847, 
    0.436938244233977, 0.717608196438022, 0.132796563375914, 
    -0.265297170155848, 0.811047089483928, 0.360597236090981, 
    0.103974644246954, 0.0566186373041369, 0.0766734366897245, 
    0.0943310173746026, 0.0628750772294632, 0.0279525471606168, 
    0.176409667340393, 0.088333944572664, 0.00490215690874474, 
    -0.163567738144123, 0.0532859229915762, 0.335204015678486, 
    0.457789361477781, 0.23716470010387, -0.136149011841875, 
    0.292671621736732, 0.345921160344096, 0.178718463614599, 
    0.286903690567043, -0.438841245167104, 0.523501548678651, 
    0.50326890333327, 0.0677599197637307, 0.0753242217211674, 
    -0.40672424655903, 0.587564296874991, 0.54587913976475, 
    0.162323578354984, -0.0425463059640799, 0.0943283849850813, 
    0.435727101927001, 0.110632893331369, -0.0809436923274672, 
    -0.0219343015482193, 0.295969713429963, 0.252885503732617, 
    0.0273118990776272, -0.0914406880434595, -0.0867965938024935, 
    0.240203427633333, 0.146503253217475, 0.077581166702979, 
    0.17752405989874, 0.138122693679686, -0.126960393042533, 
    0.0479164105508613, 0.266112054955242, 0.157144800024576, 
    0.145550887450864, 0.160675707379434, 0.0502835852838637, 
    -0.000405039086857129, 0.0170474052152203, 0.0797678445244965, 
    0.0635678447314263, 0.124022694920722, 0.0158083605055775, 
    -0.0637421491431834, -0.0325494548464025, -0.103932286458016, 
    -0.106471265189404, 0.0265233386305793, -0.0293540917625782, 
    0.0506219018391052, -0.0983140715416688, 0.0191587238279894, 
    -0.0596502457604872, 0.0300416821092263, -0.126917374115032, 
    0.0144001832048567, 0.064177474644605, 0.0685550446349533, 
    0.11643940666537, 0.15627811449176, 0.108587744800303, 0.110406886823022, 
    0.244844332343975, 0.115523430787233, -0.11670824320398, 
    -0.0186071387280808, 0.474914407480184, 0.337724422467354, 
    0.0502873674601484, -0.107508762209848, -0.19937157437271, 
    0.587797265286719, 0.266689322847203, 0.135327486131026, 
    -0.145665199876531, 0.0829855644479704, 0.235612849273398, 
    0.438982942949859, 0.403948330002337, 0.169693814640181, 
    -0.342881161853886, 0.536295944452216, 0.158011038212039, 
    -0.427404573625168, 0.0522796303778377, -0.354857715005329, 
    -0.0998340437848333, -0.284069534331339, -0.128236144102433, 
    -0.251996927671085, 0.00467382665530965, -0.300045349937292, 
    0.0121579823194431, -0.282147391183988, -0.0885489843568625, 
    -0.0628731621733171, 0.0649511188742318, 0.050155938097085, 
    0.0685562086124048, -0.0767900776308327, 0.0390744008791941, 
    0.0119249885656774, 0.0545194049415902, 0.0390956204015102, 
    -0.0694955304985845, 0.0120769869318271, 0.0540262709266771, 
    0.0569748351512411, 0.0888154931418709, 0.104456946273488, 
    0.0557024188357627, 0.0817466054287536, 0.15948759554888, 
    0.0894555327590284, 0.114093491333683, 0.18147991115742, 
    0.0179620167619453, -0.0706367565111946, -0.0780005132002851, 
    0.559956741434245, 0.448425303382019, 0.149827752423626, 
    0.0252627621015687, 0.592674146746049, 0.325343731815342, 
    -0.252634534306924, 0.522951782440514, 0.454465087747519, 
    -0.278048114488133, 0.0943088664548818, -0.552695019764195, 
    0.653870615228699, 0.324064644515266, 0.0531243874570732, 
    0.37454774824109, 0.376217127061245, 0.164477772939931, 
    0.084826459037993, 0.0843558817667607, 0.0930916571401809, 
    0.0692815535731504, 0.064134123066362, 0.0886512255453667, 
    0.0236561710272528, 0.129048715205536, 0.321964468964114, 
    0.120959833518227, 0.0727421997944748, 0.247570521420275, 
    -0.00855276880309003, 0.714980778788824, 0.448012552186448, 
    0.0139474949588897, 0.0304964271040543, -0.100690495697163, 
    0.0678024767567808, 0.91089303668651, 0.509918252498081, 
    0.316483210462342, -0.463068898995956, 0.184840123193011, 
    0.509713915267188, 0.134661705916823, 0.891522600011488, 
    0.865158333594018, 0.291993986776713, 0.253761845314489, 
    0.116815838996211, -0.149650388584087, -0.389957241763032, 
    -0.105450985458696, 0.205146792449451, 0.0468887200139899, 
    0.104937827391605, 0.19939355450698, -0.120386527570497, 
    -0.113575528137591, 0.0272048565491695, -0.158011958288057, 
    0.0572531699876255, 0.0176845622983011, 0.0658116403097995, 
    0.0839114828141871, 0.0432905677272364, 0.0503221967410249, 
    -0.0329415260619096, -0.0169598725816592, -0.0467286086441175, 
    -0.00737432788535249, -0.0473730247157773, -0.0542221382207359, 
    -0.00394132064487704, -0.0529096753062191, 0.00855523530160075, 
    -0.0523738628431405, 0.0264498133507751, 0.0543852963756369, 
    0.0822397833230142, 0.11433356172943, 0.165771909094893, 
    0.151692781059725, 0.0807256519075373, 0.0747084318622073, 
    0.222173121490603, 0.127675037568652, -0.0541234620286685, 
    0.147798674038907, 0.638197600063964, 0.160631549281862, 
    0.105618868953458, 0.0638590058408557, 0.418760607157873, 
    -0.096953350477746, 0.260730783877483, 0.826654299312067, 
    0.146365510878994, 0.0155691314112628, -0.000680889540616403, 
    0.0108427007997531, 0.0283479489814366, 0.00843844872156221, 
    -0.010670267180495, 0.0104657201556429, 0.0300081239382861, 
    -0.00704524225444966, -0.0204300151779888, 0.0496879752037698, 
    -0.0457683771010477, 0.0385670405748948, 0.00109342666022093, 
    0.0568062314266508, -0.0643090488037256, 0.0415924576476364, 
    -0.0841047226954067, -0.0260597263972882,
  0.342477901555564, 0.4771078606805, 0.294638288498854, -0.389223754018356, 
    0.27862993670177, 0.497041612983116, 0.139157399874404, 
    0.687532665742767, 0.508585130045314, -0.203798934824659, 
    -0.192859906402482, -0.0440968186831604, 0.211352602772877, 
    -0.0136976178350012, -0.162009559368512, 0.177284192265701, 
    0.169730001596454, -0.059488866391445, 0.206994270132429, 
    0.111542832107057, -0.337899294409942, 0.207080029251755, 
    -0.74384434612113, -0.276472698523234, -0.176545122612137, 
    -0.43732577397629, -0.149330148317486, -0.324319802097463, 
    -0.133558053954904, -0.260353463535099, -0.0478708239694482, 
    0.0988850412096401, 0.0745734926029951, 0.0596995385626482, 
    0.0800174444481969, 0.108913494807847, 0.195625664027212, 
    0.127813946272758, 0.00602939364436378, 0.0868248477422559, 
    -0.0594583929726512, -0.0185227433291971, -0.0268389030944792, 
    -0.0178779073988308, -0.0248021327722912, 0.013588339640915, 
    -0.0166965035497951, 0.0395018170465322, 0.00451839335873236, 
    -0.155644722317088, 0.32088281470524, 0.210711584650338, 
    -0.0576214531061035, -0.347378732301056, 0.0904551907630906, 
    0.692957775639382, 0.26261889345192, -0.157454524360511, 
    0.274667654599426, 0.451462815565402, 0.111066483728693, 
    0.163516175930948, -0.237182183273856, 0.713303020499, 0.773357056036788, 
    -0.0185089900978603, -0.00514787433851698, -0.293330325535795, 
    0.0460923621562612, 0.484104094617322, -0.160999792394372, 
    0.0020268722083026, -0.0472445414947209, -0.0316263704563226, 
    -0.0389672459999325, -0.00752006736106589, -0.0494240372871744, 
    -0.0188997515589474, 0.0354750973844031, -0.221060757869294, 
    0.0115330732912787, 0.456824337932354, 0.0516271886197996, 
    -0.155159286725775, 0.149975169200416, 0.274112301348633, 
    0.212918660267047, 0.808959189596788, 0.670111230847248, 
    0.11837075161808, -0.0740729529958578, -0.0724614776144159, 
    0.171659357273365, 0.258818138389872, 0.188244130192543, 
    0.098905485852215, 0.0437365888054057, 0.185693459994941, 
    0.166546565861842, 0.0214894000340093, -0.0642707798553581, 
    -0.0793492061724055, 0.0204251854930881, -0.0853085830780361, 
    0.00282494306908093, -0.0567135310786718, 0.0235982518069032, 
    -0.122324683718922, 0.0171791206204249, -0.0839009352638469, 
    0.0082119878403811, 0.0278959205235309, 0.0695316046206827, 
    0.0566523036768538, 0.0248566022436319, 0.0476639369881521, 
    0.0896349103612375, 0.0322761621069267, 0.0102204857024191, 
    0.149188071538889, 0.384699876534362, -0.213095789377974, 
    -0.327151346460785, -0.372513405856173, 0.723565979676568, 
    0.481305836379089, 0.142890362203556, -0.00640516766052189, 
    0.231924531701478, 0.232374818217403, -0.149150059626413, 
    -0.160235002983488, 0.520888080086885, 0.288927490087378, 
    0.699485457614963, 0.7862894377722, 0.0653165982548082, 
    -0.0470687664848064, 0.113159134814127, 0.626489991325866, 
    -0.0460508696584945, -0.0200382900041141, -0.0639304299044871, 
    0.138858256247181, 0.168969076412481, 0.174433084372054, 
    0.132586738680788, 0.0429116307810153, 0.234940891291318, 
    0.142481066916046, -0.0551504474375461, 0.531055098484637, 
    0.355249419096586, 0.14644439426868, 0.463517923919485, 
    0.247039934276685, -0.0547089879699312, -0.12901683677369, 
    0.0741236773500552, 0.386692894257702, -0.0580321898122258, 
    0.000167671088537283, -0.0529428223642622, 0.00114977072506807, 
    -0.11649473108046, -0.0697100969115854, -0.0650881768275315, 
    -0.0732144320756804, -0.0606318107208042, -0.112930238276214, 
    0.0821720520089574, -0.110368683862629, 0.0665886930637999, 
    -0.0711547039994352, 0.0459145051979337, -0.027228827862078, 
    0.0778450694975445, -0.0456414520771317, 0.046641952093494, 
    -0.142490529045443, -0.0267418374962248, 0.0565068558249541, 
    0.134380179369858, 0.0842950728657432, -0.0425326070187041, 
    0.160839062824309, 0.22390724308797, 0.0169796330682693, 
    -0.0250904506477083, 0.0749488378352081, -0.0660302834193131, 
    0.405026049805718, -0.222139554735477, 0.302492523723899, 
    1.01349853691294, 0.067558119651091, -0.194086301939859, 
    0.319700448260618, 0.456730472361654, 0.0921137100991095, 
    0.118082485100979, -0.16609736326886, 0.461224095034407, 
    0.34313528542253, 0.222129764241013, -0.0799406365879466, 
    0.207977373817923, 0.388225033202979, 0.303338761261358, 
    -0.0829783963127714, -0.395353304751607, -0.104785721703311, 
    -0.242557331414062, -0.144118164434325, -0.14913600201629, 
    -0.23164817688172, -0.0476956187362461, -0.164094719860006, 
    0.0144834261080884, -0.178681221909392, 0.0727071723780947, 
    -0.0188220942665367, 0.0850101155303324, -0.0282831857093094, 
    0.0592037261801574, -0.133234662366282, 0.00255963676300114, 
    -0.0831951434350542, -0.0929446131830453, 0.0338137537399414, 
    -0.0206196125750953, -0.01104569874913, 0.105792851959075, 
    0.0920821364609632, 0.00535645435019147, 0.218023443655157, 
    0.219314384241734, -0.115953515365277, -0.053302138026146, 
    -0.192989403936986, -0.134742390361469, -0.16803282136694, 
    1.07250359056627, 0.0978670043962625, -0.161004612321098, 
    -0.296981598657285, 0.362996509563534, 0.53287334651982, 
    0.512065378012465, 0.4668849326348, 0.0411234678224248, 
    -0.201502178943776, -0.11609863968436, -0.174130641431998, 
    -3.73137943176505e-05, -0.199799426066257, -0.0733320155755898, 
    0.00155575059161761, -0.122638040572849, 0.053350483395971, 
    -0.140761348416844, 0.00562816038539997, -0.109157443677543, 
    -0.154379635653347, 0.170036484409057, -0.0307747105158568, 
    0.112003779526232, -0.203279294714002, 0.00664205599455706, 
    -0.0736624324193633, 0.0117817987684334, 0.0824883960269712, 
    0.0217656855550565, 0.0339729694270323, 0.061100318169799, 
    0.0446390374332343, 0.0744108355308319, 0.0897394947753185, 
    0.0918506369850121, 0.0564376088515285, 0.0695518743574157, 
    0.0520530386313501, 0.0684331342813813, 0.0651177384348282, 
    0.0771392638889647, 0.055918467965856, 0.064227594977709, 
    0.0597798512652163, 0.0656382194931405, 0.0373698376504914, 
    0.113368442334792, 0.0508420615146846, 0.0866273084019061, 
    0.308219228116475, 0.182607400019729, 0.00618567108017007, 
    0.236798207633292, 0.272551118587687, -0.0202321923513753, 
    -0.00691714707437605, -0.0380128535540998, 0.611832392173697, 
    0.00631796654951648, 0.531982935406985, 0.80942632038091, 
    -0.0997013665231973, -0.0792836621858187, -0.0937371673268084, 
    0.851521717383628, 0.250011995265316, 0.179924698533878, 
    -0.281719123762848, 0.140025673968229, 0.282947592637679, 
    0.436374290916599, 0.310718724288738, -0.0246617683436649, 
    0.108562183981168, 0.728973485747836, -0.105048708473079, 
    -0.141362567880416, -0.0650435275752129, -0.111528146807427, 
    -0.106738540532739, 0.0314283435601111, -0.132356232326799, 
    -0.0200353309973765, -0.122642833239939, 0.0145987786526261, 
    -0.0617771961449173, 0.0968001141426494, 0.031338760133911, 
    0.0531445802189988, 0.146457742301803, 0.102439470033147, 
    0.0478226037536911, 0.129808254450377, 0.128523376935014, 
    0.0623192803777085, 0.0480582925386432, -0.0274124948561828, 
    -0.0416920947478562, 0.015574573844032, 0.0301634982639626, 
    0.0499855778455955, -0.0236959571189318, 0.0419768053431319, 
    0.00113189535596232, 0.0505220080757395, -0.0550941393619529, 
    0.0514313560560371, 0.124763719636275, 0.0321568128561327, 
    0.136075705340355, 0.265816859216056, 0.145441717023057, 
    0.0638300363059188, -0.0872742626022674, 0.102887287700238, 
    0.210878658394757,
  0.116689422978001, 0.123735570278537, 0.121201059726097, 0.117050184645422, 
    0.118501818152037, 0.122994122498095, 0.13771722348079, 0.1434516702855, 
    0.106602746915485, 0.0709375246433716, 0.138967087477404, 
    0.149896228769894, 0.100020257194319, 0.182619506461803, 
    0.280223975686204, 0.208279618410933, 0.15489193154662, 0.12594540617479, 
    0.0883023746614457, 0.477626234500359, 0.328749507746391, 
    0.0495909135291329, -0.120773668109813, 0.549386302581841, 
    0.333826697197276, 0.064549413765885, -0.12257084292761, 
    -0.100689091420149, 0.62713229425619, 0.0917585350111406, 
    -0.0788505468295028, 0.026880450072357, 0.103701903367911, 
    0.12300769724264, 0.587260374553774, 0.198974926117881, 
    -0.179965479894975, 0.220084211266471, 0.404918274387594, 
    -0.0468050223617107, -0.0798185568266511, -0.202316291659506, 
    0.017187649628734, -0.0619500199681279, 0.0281256654647099, 
    -0.087242527328464, 0.0410536530102408, -0.0601265958682121, 
    0.0416442947880895, -0.19126059459878, -0.0398593251377591, 
    0.142349527378018, 0.201307970942217, 0.140952457552892, 
    0.0518646524851426, 0.196085683213063, 0.473387140782508, 
    0.24113122539995, 0.00996253700759658, -0.039713245580456, 
    0.797473304401673, 0.12988497883164, -0.342005680554299, 
    0.22991578924387, 0.642971872215373, 0.0288036022874606, 
    0.120228972059777, -0.282741218063833, 0.529716531113636, 
    0.351355698664859, 0.148762719064586, 0.179410047372994, 
    0.0692093280652242, -0.245105911365482, 0.229755149335547, 
    0.523190117405594, 0.194958433482016, 0.180412352388614, 
    0.618843301128869, 0.194517107036358, 0.0526244519436784, 
    0.141881112521099, -0.0385824564804973, 0.198346657347583, 
    -0.0356384228984339, -0.151532124237284, -0.229159634059264, 
    0.0404068054547159, 0.0184915608760446, -0.108139340920196, 
    -0.0503116508298575, -0.112537316023797, 0.115903719173775, 
    -0.113552859616313, 0.086309491652604, -0.235421789521431, 
    0.00826881875522134, -0.154914288718517, -0.00197285768024977, 
    -0.263225875073736, -0.0599183440538331, 0.0833411389648386, 
    0.110583212146002, 0.0746342789438406, 0.137944306593268, 
    0.233469727712253, 0.245615146750745, 0.226606484187767, 
    0.166551819750398, 0.0837693360987393, 0.167670643431233, 
    0.337222272475392, 0.431239338082707, 0.295368802124193, 
    0.0797502062686246, 0.201436778881791, 0.689201831553394, 
    0.373478221325655, 0.0703072955213959, -0.0413301129154398, 
    0.634747471305497, 0.334493032681416, 0.07530148861461, 
    0.109894489075868, 0.390791936931768, 0.0981039817350167, 
    0.16361879841161, 0.630551639831598, 0.495328632429273, 
    0.225681323615524, -0.187277442998175, 0.280212979998926, 
    0.283961564427917, 0.22432291828313, 0.364667001757386, 
    0.228288357334435, -0.160973610640153, 0.537282208905872, 
    0.305550458188389, 0.0274099329332194, -0.0606182363893168, 
    -0.171536393000112, 0.0704400601069004, -0.124990416727606, 
    0.0190924128303598, -0.138719431130835, -0.0147644651684167, 
    -0.0179852038349723, 0.104427214497579, -0.201447509165121, 
    0.103238960533817, 0.247129226002751, 0.0998823440703509, 
    -0.241570297819987, 0.254990405837471, 0.489401674194651, 
    0.172040888126008, 0.040271195690725, -0.118448032477386, 
    -0.0267497232592545, 0.364285638134735, 0.416542795665405, 
    0.32754861923174, 0.355265445831409, 0.382838683356943, 
    0.237192419872015, 0.081209894864637, 0.336796815664297, 
    0.519472746633709, 0.201824569226401, -0.0771032535492612, 
    0.241534861444481, 0.313718185861338, 0.310953653750546, 
    0.532829013229211, 0.263109606535593, 0.0849363805912277, 
    -0.165083345431585, 0.881696016921703, 0.0169295027932165, 
    -0.247963319294652, 0.0627992193499631, 0.473637500486444, 
    0.398048676744888, 0.443802528091389, 0.133852502686674, 
    -0.502503795308696, -0.156981208825474, 0.482040266345081, 
    0.626902337900647, 0.497507364581178, 0.189286922567922, 
    -0.0409574701433935, -0.0424130156143008, -0.033218538960516, 
    -0.0929105831838909, -0.028222758854982, 0.0967582242257405, 
    -0.0313698936793846, -0.0479174812856173, -0.0150896091906392, 
    0.121544193189954, 0.127751706985985, 0.10689749422846, 
    0.162158174794736, 0.129355572265771, 0.0265168760900028, 
    0.0852135560994602, 0.184800306479718, 0.110127982106684, 
    0.0692094408640557, 0.111814112163071, 0.146352282671102, 
    0.189210010105891, 0.272292919753138, 0.220693116622691, 
    0.0988539976020216, 0.00889256467533471, 0.211123006404649, 
    0.254835629142725, 0.124291872538391, 0.0875244296743777, 
    0.104042825775027, 0.103921192060084, 0.104985576482763, 
    0.0694296910808866, 0.077376372536914, 0.102639200569534, 
    0.106718118257313, 0.0434241001125968, 0.0743887528911301, 
    0.0186996835763071, 0.441006224278378, 0.253345682845017, 
    -0.0727559269206178, 0.299282731898983, 0.462688358652214, 
    0.118331361199422, 0.0238628882324899, -0.0646930340995782, 
    0.102377553976713, -0.237306259918925, 0.941985257703083, 
    0.402298180051389, 0.0655789192598807, -0.02174399737983, 
    0.0295629580001321, 0.253615602114164, 0.980571389344958, 
    0.0433179493505856, -0.200368984744512, -0.187067026950077, 
    -0.0702581607680917, -0.0268778654859177, -0.106263485809644, 
    -0.0433083197587548, -0.146439389864364, 0.0140348218862755, 
    -0.278222951000227, -0.0152693524233134, -0.140779852867264, 
    0.0772803290633504, -0.165936366047382, 0.0107980466424924, 
    -0.155570280058726, -0.0565566351057427, -0.0673791164966241, 
    -0.0866808620740959, 0.00956864202624402, -0.111929612064699, 
    -0.0484033256877867, 0.0757509379178074, 0.124716882372195, 
    0.107382475676811, 0.0939999712803294, 0.0936140962955846, 
    0.111798422061242, 0.166212505704266, 0.135783114921455, 
    0.050226004464953, -0.0050019869290221, 0.269008811153741, 
    0.33449111743479, 0.12305696302734, -0.0183349468859904, 
    0.316826756932133, 0.463484047895983, 0.359737753411746, 
    0.160743565864475, -0.304281587315811, 0.19013604088857, 
    0.650056904591379, 0.0266465657267441, 0.027451435934231, 
    -0.257351034149769, 0.17502974011381, 0.407709782419618, 
    0.176006244338197, 0.406119138221575, 0.515083830597803, 
    -0.0599675277414221, -0.0750906701097496, 0.0187350143557326, 
    0.0877680316188728, -0.0530643567332758, -0.0441269606219088, 
    -0.0659576124641934, -0.0302008486892128, 0.00711166928064025, 
    -0.0578923384458164, 0.0174884535866316, -0.0552669375537155, 
    0.0379037751167677, -0.032417279879899, 0.0209675844945487, 
    -0.0320822648840522, 0.0130030292311764, -0.09259025067146, 
    -0.0273420060343477, 0.0180727247612086, -0.0285579868832259, 
    0.102299677038916, 0.165537905830608, 0.0850018307673394, 
    -0.0102829519894935, 0.180169125349707, 0.146529671352579, 
    0.0215571416499746, 0.0891307519554168, 0.305761546450614, 
    0.402243407178401, 0.0589859150341272, -0.0236301502352689, 
    -0.463053660358339, 1.05464619441261, 0.55061396900838, 
    -0.17447525971051, 0.855597323887919, 0.542891346600525, 
    0.0339818349651252, -0.148292939527061, -0.0748572271512201, 
    -0.0869325636733737, -0.124180435122134, -0.0355450790851184, 
    -0.124121718575351, -0.0634598451521793, -0.0783687501421545, 
    -0.0411825920058051, -0.088373946000338, 0.0194508238666522, 
    0.10040894367825, 0.131354816369129, 0.153580806616565, 
    0.137116079624705, 0.145368930086955, 0.184099819021726, 
    0.17583169542596, 0.135529524720518, 0.131515059239836,
  0.339280820309065, 0.282884987285653, 0.19594648036245, 0.113149356061336, 
    0.030028576235041, 0.0211312347802898, 0.362211386265934, 
    0.407585955665551, 0.229429637996276, 0.116682842360854, 
    -0.266971740623192, 0.104088991437168, 0.483807086655919, 
    0.346559844170273, 0.110678353541044, -0.16602716682573, 
    -0.116500820505716, 0.348527224208756, 0.4469857530957, 
    0.230125483336709, 0.0149685595670462, -0.0350812077516061, 
    -0.0514157303920103, 0.389439868311201, 0.361232799880197, 
    0.129269843249074, -0.0360267934776935, 0.422783236192343, 
    0.107013010266814, -0.0287470248076003, -0.126278296629615, 
    -0.0894018161477978, -0.0270024376756759, -0.115734376496856, 
    -0.0218345558299729, -0.142635734146926, -0.0561729620351422, 
    -0.0820509245580661, -0.0382989943648432, -0.104574266546924, 
    0.0910889198866867, 0.0888040873917644, -0.0309930753311038, 
    0.290468114063128, 0.234514649081635, 0.0453852301309042, 
    0.0102349177175133, 0.280576858500291, 0.389055764868089, 
    0.200685646754585, 0.34991331137296, 0.405218340550024, 
    0.293944445032344, 0.801048141334245, -0.0131318893798018, 
    -0.290779846935674, 0.573747699809702, 0.0804012271125718, 
    0.823135174435876, -0.0363510565592936, -0.143491826405384, 
    0.0411287739418175, -0.353361653822284, -0.0677361873646266, 
    -0.16567787079427, -0.227421963877897, 0.086608691312629, 
    -0.186882171803138, 0.120564476361965, -0.254296903573285, 
    0.0180307110169743, 0.0955777725118952, 0.121150508295287, 
    0.110987537178025, 0.144915200789304, 0.132790347014068, 
    0.154939575430722, 0.172463040964603, 0.175508368738319, 
    0.106926991504981, 0.109396447220349, 0.13642175032913, 
    0.148026951044871, 0.145178356446507, 0.190848718820326, 
    0.250582374074441, 0.210348874979018, 0.14111754978733, 0.17883775447948, 
    0.265197814049644, 0.214941511481294, 0.157307655655825, 
    0.136643799923252, 0.153961865268059, 0.16482442751442, 
    0.135429314177418, 0.126601204924015, 0.162779198162576, 
    0.142894366559541, 0.106821247968594, 0.199252690457795, 
    0.173165836160305, 0.0838837521093434, 0.299304095097569, 
    0.302000920980907, 0.0794271649191616, 0.0909493093836684, 
    0.376589483985709, 0.261912529469067, 0.35683706667382, 
    0.277100853381985, -0.190927017980478, 0.0933026159630217, 
    0.492993820729067, 0.294514416676897, 0.0858415630183436, 
    -0.185949049675032, -0.102875999153693, 0.510180702900729, 
    0.31009991362107, 0.0276193808980692, -0.00309548739700137, 
    0.290065904743366, 0.1030185279275, -0.0622480513435756, 
    -0.014032565715979, -0.135378189429264, -0.0791192680155527, 
    0.149811465961871, 0.143860666940385, -0.116222835182526, 
    -0.135131705455132, -0.29306572867421, -0.113260502719614, 
    -0.112155838409931, -0.336761057604287, 0.121499872413316, 
    -0.0788792517883568, 0.0410388348690951, -0.288544072316303, 
    -0.0452231829153386, 0.0458995291816128, 0.119517209063541, 
    0.128393581884711, 0.129559657607989, 0.110927139598233, 
    0.126157940248858, 0.19750764955041, 0.171760818633866, 
    0.0991452336800576, 0.128884481650419, 0.153529489498061, 
    0.264418257570696, 0.371510838886182, 0.219315200074105, 
    0.0295551054717417, 0.492860107424426, 0.297937885848962, 
    -0.106648138834471, 0.328224380067239, 0.507716011635901, 
    -0.178211919886302, 0.0670953748421574, -0.367754374895693, 
    0.517692275037876, 0.363489322134486, 0.155902578833054, 
    0.0833201018133186, -0.213510961678513, 0.327886900159119, 
    0.359140525966824, 0.0906711734332039, -0.0340466565636025, 
    -0.0455265113044915, -0.0256442015464417, -0.0600799329930456, 
    -0.0806816481020974, -0.00664872781047948, -0.078296694390292, 
    -0.0857078603335584, 0.0308601834404741, -0.0834874763672627, 
    0.0756315970147406, -0.0881917158372076, 0.0196835954479558, 
    -0.104234187914109, -0.0430975050221136, 0.0174572659919513, 
    0.0192150948711761, -0.0941449925041554, -0.159152068751603, 
    0.0718384195753835, 0.300595270165023, 0.109073445067311, 
    0.0387385115736878, 0.0629093828302818, -0.193750893656317, 
    0.265126607733748, 0.341795964134254, 0.13145319502443, 
    -0.0317052296718982, 0.0410867782665649, 0.410743089532612, 
    -0.197858130966656, 0.391219311057963, 1.2270552928088, 
    0.0139990732447841, -0.392328378984184, 0.365050603946992, 
    0.511949031431043, -0.156603883351364, -0.0889271797093024, 
    -0.105316502763907, 0.0165946017445159, 0.461463948470026, 
    0.192809143631516, -0.0863232497849263, 0.1704831099755, 
    0.315803777144011, 0.0111608322835597, -0.0871785079912742, 
    0.00705775278674986, -0.13759348288979, 0.269334918860375, 
    0.0269616720706171, -0.100708007691803, 0.0243123654408059, 
    0.120102112416095, 0.10955088776046, 0.148998032712334, 
    0.0381216594403754, -0.0404595075773217, -0.0148031783820293, 
    -0.0724236786757907, 0.0277526017583319, -0.00470887301344448, 
    -0.103051035331349, -0.00249307013998717, -0.0543212745532129, 
    -0.0576860227982504, -0.231993549365553, -0.205274220089431, 
    0.00841482134742395, 0.0870958215061428, -0.520464709191632, 
    0.174435116318838, -0.263062039921471, -0.184291060402275, 
    -0.0377966197528324, -0.478125642189928, -0.125292599879316, 
    0.0200687523248905, 0.0135706514760559, -0.0299775904254985, 
    0.0356538544511812, 0.0706663062716013, 0.0797159092952008, 
    0.121540168969581, 0.107743834084297, 0.0674204007631572, 
    -0.223419510828056, 0.020703904588517, 0.608721517150163, 
    0.129063507707541, -0.324633461039373, 0.245452617571713, 
    0.525808896674092, 0.0017862844078909, 0.0634244036045732, 
    -0.333838177472973, 0.431342679143377, 0.391437913696543, 
    0.162925454718324, 0.188563354268409, 0.357749378579857, 
    -0.262165814130029, 0.580343875433604, 0.420197653124722, 
    0.11558807648417, 0.0848209899226859, -0.0496319401856148, 
    0.332305868629373, -0.139501651597497, -0.0947392066169676, 
    -0.0696994344934333, -0.114873240271532, -0.254507406528982, 
    -0.267100419295659, -0.0161820872324147, -0.00948654307009816, 
    0.103170977787729, -0.183612055357533, 0.0485393985385382, 
    -0.00651164169154735, 0.0349908788618323, -0.314076200815548, 
    0.0368909146319131, -0.148366158011362, 0.0376711204102993, 
    -0.382897033138247, -0.0424418851573714, 0.0404748854042051, 
    0.0669542655667763, 0.0862484500165095, 0.110759136775158, 
    0.118721248898608, 0.092325129981309, 0.0100369765177487, 
    0.0541883814051943, 0.00251871351952926, 0.107298936689686, 
    0.127717751330345, 0.143640854980248, 0.126995464174651, 
    0.151086856510167, 0.104263402537234, 0.321501929878172, 
    0.317912858154357, 0.0277300001069486, -0.129382824199885, 
    0.404525770181594, 0.330076184234139, -0.357940519512328, 
    0.335948362820838, 0.462846169601803, 0.440513855567463, 
    0.818501658635178, 0.29016391730118, -0.464148512720561, 
    0.178870299664213, 0.801901596060851, 0.0796639932177816, 
    -0.23072433174751, 0.0996444236822933, 0.374523074713625, 
    0.552867154893705, 0.349387864156245, -0.151150323198072, 
    0.415345326659286, 0.731508957751494, -0.14574388045557, 
    -0.158471562961883, 0.127126501366403, 0.0868141839799871, 
    -0.0819675458605464, -0.0100687374887926, 0.182114598104581, 
    -0.0387664487158462, -0.0351260642626096, -0.0792458009480624, 
    -0.14126395400257, 0.291587815792789, 0.162138379425642, 
    0.0724097116104157, -0.0375038723507198, 0.276027828347182, 
    0.157563709152882, 0.0130989227721429, -0.041233321705608, 
    0.181674653763306,
  -0.225909219653459, 0.111126876535562, -0.169827377010899, 
    0.0410444725328471, -0.445791221060505, -0.0566513551593582, 
    -0.115700511941946, -0.163323120653378, 0.111965729841973, 
    -0.355705430674489, 0.020754784277032, 0.0800083631889092, 
    0.092061904623148, 0.136754361027763, 0.23442408097715, 
    0.263208098005535, 0.265508648469215, 0.292997124128367, 
    0.251422675182467, 0.201956864743662, 0.327717531609439, 
    0.359695530596677, 0.261718688078821, 0.323000650390088, 
    0.493724054887017, 0.317495762155222, 0.109636843651038, 
    0.501879682468544, 0.575463276764109, 0.197647092007218, 
    0.0652964526583159, 0.624432611688375, 0.409622676187802, 
    0.10628727018874, -0.212999495097969, 0.19644324496936, 
    0.554463283249981, 0.11751725850861, -0.140446995834583, 
    -0.0536979542320706, 0.418227939536595, 0.417302743936529, 
    0.194970464848994, -0.225948684821805, 0.217803575867686, 
    0.434862860711523, 0.198237011123815, 0.0715795520081882, 
    -0.00764612216792276, -0.110449968422274, 0.538553410226844, 
    0.280456902285933, 0.0281884279918931, -0.191042381358928, 
    0.09154245894358, 0.530281146228051, 0.127212431048893, 
    0.00338433397849744, -0.0766568029476392, 0.119032203637254, 
    0.247796906735522, 0.246790586655586, 0.0203471385173023, 
    -0.061932205773043, -0.0226410726568931, 0.0758777428467481, 
    -0.0586192554599724, 2.28613394386845e-05, -0.173978310010201, 
    -0.166286983220707, -0.0395146750595738, -0.0823635420008961, 
    -0.0461949570742593, -0.101606770180191, -0.0271041939041775, 
    -0.0837449351297605, -0.0157129023459319, -0.0670947254888184, 
    0.0411962717784611, -0.0853562982989685, 0.0423890199190111, 
    0.0539018724439359, 0.0646662811608536, 0.0656572495654445, 
    0.0721748669944053, 0.0529569783383974, 0.0400245244455411, 
    0.0817746400716644, 0.0576122155916927, 0.031385040322227, 
    0.282432049037856, 0.165714672657123, -0.0838936954212261, 
    0.289787620047435, 0.369411496158677, 0.210657657093304, 
    0.173109800883446, 0.261452534723311, 0.224436680454167, 
    -0.23700258195429, 0.707164472916661, 0.444341180565525, 
    0.174045110710282, 0.0874716271932442, -0.140347597634463, 
    0.107406094942577, 1.17074176509424, 0.117103656380609, 
    -0.0142291258680964, 0.128120685726113, 0.0134962167820499, 
    -0.193626302276285, 0.237712106408068, -0.153661203644078, 
    0.172504665578912, -0.0943894058923197, 0.189051399489306, 
    -0.100983883802353, 0.168139029635435, -0.209382464527821, 
    0.0993248364985832, 0.148725994631562, 0.201478500938859, 
    0.191762368307145, 0.186084991752048, 0.0374472301157462, 
    0.0991922477489527, 0.145235296159772, 0.075213139855781, 
    -0.0443922079364206, 0.00501780856754308, 0.00560879677411105, 
    0.00787674013030648, 0.0138930859092447, 0.0130239961945059, 
    0.00539905727082972, -0.000624491275560773, 0.070610671319685, 
    0.145350109555603, 0.0131524069165955, 0.287449521827943, 
    -0.119456854110515, 0.271598199308918, 0.598101836619593, 
    0.660311364452608, 0.270719881347675, -0.284271117622002, 
    0.103887319503074, 0.591978666246769, 0.347219156379582, 
    0.0482574951115706, -0.178833568779247, -0.247122697497162, 
    0.4043653274627, 0.394446837657099, 0.635834981181775, 0.333477094468629, 
    -0.313541572360538, 0.2073229133374, 0.615098451263432, 
    -0.222654793376086, -0.150447333258304, -0.00952657960551587, 
    0.308317232140278, 0.00888968833284008, 0.0185763291437548, 
    0.0288637657787727, -0.148575053028186, 0.243647512425197, 
    0.195225228641713, -0.0541131953722814, 0.304375148691009, 
    0.385370584940607, 0.122827693849327, 0.0551170605286053, 
    -0.0371094156744932, -0.247177235831052, 0.291967567953651, 
    0.298531956604986, 0.127713100324371, 0.172542118485481, 
    0.254427338538984, 0.113003011048098, 0.117829958754745, 
    0.302490520139978, 0.102088294223306, -0.00903581670490858, 
    0.0828659510208752, 0.219846551711163, 0.0854105885050479, 
    -0.0124952739201697, -0.0498655406331612, 0.0397986616805506, 
    -0.0183905181748797, 0.0379910216327843, -0.0203553098390349, 
    0.00781123087961372, 0.116728430264599, 0.124733716643246, 
    -0.152690977061838, -0.101319123168117, 0.273110922209689, 
    0.400989188986655, 0.1580000278843, -0.0996881730810559, 
    -0.0777628389481221, 0.309714239339833, 0.626330411841693, 
    -0.0767439543373417, -0.148764269734993, -0.423379466102663, 
    -0.0633682660055756, 1.03485386811843, 0.0299629248564648, 
    -0.381244170092079, 0.0516462114351014, 0.686618760093475, 
    0.181516543440154, -0.0461090812624795, 0.332070290334197, 
    0.548951637662783, 0.630620270324514, 0.327874634268596, 
    0.164980808759868, 0.57272975770776, 0.264769639258379, 
    -0.0278005357938336, 0.320927579847944, 0.268378790206021, 
    -0.0778510494223687, -0.0775116835142125, -0.097098536603853, 
    -0.000840068197506025, -0.0781728762510389, 0.133087068762906, 
    -0.0795187950774993, 0.144749580483804, 0.207632487879702, 
    -0.150274509536711, -0.0639357944798053, -0.0475551045945768, 
    0.00143821782205304, -0.0125346025834528, -0.00196509001410522, 
    -0.0193877025524115, -0.071238642299122, -0.0344920608468184, 
    -0.000151193907629521, 0.0713920700633573, -0.0633215974047202, 
    0.0256447315063208, 0.055546992371146, 0.0567958487039262, 
    0.0564757886253515, 0.0633300786409295, 0.060610495251666, 
    0.0456484293188126, 0.0794078518671296, -0.0487858792801279, 
    0.0950753624336967, 0.459268409853784, 0.0195294893883323, 
    0.225068700246116, 0.721117185864612, 0.221652660300995, 
    0.157534667670919, -0.243115420756658, 0.0548133577161048, 
    0.30273020985204, 0.333851650999099, 0.497866690018742, 
    0.378368762904437, 0.12031795367222, 0.175766245893348, 
    0.379003450232366, 0.0639821088504807, -0.0567525743195721, 
    0.10719292991619, 0.24368505803774, -0.0136162650805314, 
    -0.0574857544880608, -0.16889705527737, 0.0703252330343388, 
    -0.109963688373034, 0.0443661751203612, -0.16938262686157, 
    0.0156496248713819, -0.0847692803449535, 0.0414193070409382, 
    -0.216939243050942, -0.00723416576510388, 0.0727423043774406, 
    0.025980494665055, 0.233939046303901, 0.119335179253248, 
    0.0479674175145468, -0.070485904744628, 0.32626802093888, 
    0.0589425210234, -0.193166140545665, 0.244534996153927, 
    -0.35433655322252, 0.517798705494023, 0.867273844891441, 
    0.340370554298082, -0.0200132322284722, 0.21844086027097, 
    1.2200480572101, 0.292772873402147, 0.144179881046853, 
    -0.0224472153748249, 0.470276947563573, -0.245778278209037, 
    -0.043013279691509, 0.120556540304921, 0.185343978807344, 
    0.145065225303497, 0.186726887382153, 0.113904689292453, 
    -0.109851290784941, -0.40269684967595, 0.369442068344433, 
    -0.335547659453276, 0.170401124361553, -0.505106466273915, 
    -0.0389616266666587, -0.34890775159719, -0.267058773777821, 
    -0.0727214200739157, -0.294954902110474, -0.0147383893284375, 
    0.0420322003901739, 0.0487458703955277, 0.053988690622698, 
    0.057923468641558, 0.0405576948557408, 0.0433866976835396, 
    0.0864764981254294, 0.0455313299181344, -0.0247080222061189, 
    0.157728113099603, 0.17971060473119, 0.123271791424973, 
    0.533675915066862, 0.319354135575505, 0.0706778514083939, 
    -0.301216673944703, 0.735292623447892, 0.342207983012457, 
    0.0592561382832684, 0.216085980370244, 0.444765073705654, 
    0.263769232203185, 0.34725231456302, 0.689584936554689, 
    -0.112988295432776, -0.247685270354879, 0.167912402156648, 
    0.353177670714117, -0.0744341736413677,
  -0.431212623829752, -0.258994828760103, 0.552145726847786, 
    0.396658885416853, 0.269690096066709, 0.251519908130357, 
    0.0141232831560565, 0.150949648728403, 0.893421925583141, 
    0.0502431967224103, -0.110790828143725, -0.0245661163985978, 
    -0.0625730693352898, -0.0366840858374544, -0.0622893213793431, 
    -0.0389899043323215, -0.0457201870463326, 0.0122338497169967, 
    0.171614023578585, -0.190478913299807, 0.225656272694081, 
    0.252982914988424, -0.00753615017069054, -0.0443633505254588, 
    0.4619874539506, 0.22330559958682, 0.012038046731292, 0.156782962231425, 
    0.355046410782587, 0.380030218083053, 0.179866532290536, 
    -0.206276339775105, -0.294899699009425, 0.687581566677629, 
    0.127160489448442, -0.0437285143913676, 0.248195071922182, 
    0.4486672499049, -0.152054781419602, 0.271623147982257, 
    0.717008392734386, 0.159342289659119, -0.0427508854416718, 
    -0.114235003218893, -0.0396337571043034, 0.131900003371621, 
    -0.018286449004008, 0.198888458525573, 0.148028615967678, 
    -0.102697376857393, -0.0516732780852858, -0.116638201280607, 
    -0.00282318485001086, -0.121380236011198, -0.0743131358514039, 
    -0.0848270839314072, -0.0859823127432963, -0.0695482498839888, 
    -0.126394613370254, 0.0398977473181297, -0.0587182206359762, 
    0.0465943901181015, -0.0102779717424413, 0.0550636452458409, 
    -0.078853373415753, 0.0401303952911502, -0.0828023148168045, 
    -0.0120193597550616, -0.0395289288002977, -0.0116305046728016, 
    0.0014036662776659, 0.0457948413069229, -0.0834303112930562, 
    0.0203800487827849, -0.0204975217344782, 0.029685707827469, 
    -0.017695571715803, -0.00822524112390907, -0.167773065809677, 
    -0.0449874091671791, 0.0155578305609177, 0.0189739962124461, 
    0.0804909997324284, 0.0753253913383403, 0.0625628025807621, 
    0.0669236730117191, 0.136976307001088, 0.131277121826365, 
    -0.149677636399501, 0.162420113989161, -0.249731081988595, 
    0.358744017927352, 0.381380946728968, 0.234339768112722, 
    0.195165204709485, -0.456527767627296, 0.354156799573947, 
    0.517986016390538, 0.238110704215602, 0.0303690399456445, 
    0.198253206934375, 0.150163087914631, 0.234909550784226, 
    0.425741380849265, 0.287656145965118, 0.260314012282202, 
    0.939038347711916, 0.291913233924706, -0.260899933097551, 
    0.134327863559914, -0.283633865082278, 0.303811909395308, 
    -0.383875931330135, 0.209660324026208, -0.467510715415148, 
    0.00400534177182414, -0.388814226975433, -0.231595477242619, 
    0.12455171485106, -0.351612128307737, 0.216842011079081, 
    -0.0149900377614007, 0.0566933760836287, 0.102613361910314, 
    0.0924549383064042, -0.0175457515092022, 0.0269609830985181, 
    0.0884549939295101, 0.0868719716260045, -0.0663721275426508, 
    0.0889002251631467, 0.0583359608011298, 0.0288143791107205, 
    0.259405221462085, 0.0993654894989712, -0.0243644472614878, 
    0.083002445999999, 0.220714374946357, 0.126898599720004, 
    -0.185482673038272, 0.202842416981603, 0.724282136362859, 
    0.390116158272809, 0.200180430107589, 0.374351469546165, 
    1.10617111173794, -0.0726320136752963, 0.0076028988262201, 
    -0.135233170844997, 0.582847741378276, 0.295044152233289, 
    0.213333567437597, 0.155270349831412, -0.00829014506980331, 
    0.314045862264811, 0.160649011025294, -0.0384499327497461, 
    -0.078755879166065, 0.10320575958402, -0.125653967793715, 
    -0.267587024453475, 0.107304344658159, -0.23720091693012, 
    0.0154245739700933, -0.155806156152054, 0.0602870846316635, 
    -0.0953117867265795, 0.0814254977370162, -0.25531951913934, 
    -0.0426033527639881, -0.0353603561933127, -0.00668337923614069, 
    0.0480792292968272, -0.016106279559309, 0.0526982135635406, 
    -0.00221973353392658, 0.0478349224167586, 0.0177657610726048, 
    0.0674015459884612, 0.00701319005247568, 0.0435555791423559, 
    0.0237999628040096, 0.0377761760902307, 0.0153977720388653, 
    0.0346253435761105, -0.00295273670444726, 0.0201134355371092, 
    0.0240847790977522, 0.0111342076253898, 0.0387665710629166, 
    0.117823332262799, -0.00289753608472851, 0.219139299869505, 
    0.251464398928387, 0.112463369700774, 0.00664370503700569, 
    0.200910169793332, 0.338440595470298, -0.178479128152331, 
    0.147268061727141, 0.819510449207541, 0.106595367660476, 
    -0.342759879140606, 0.421238885505616, 0.993414680201653, 
    -0.0190437436350748, -0.180910791904518, -0.311856652404947, 
    0.366826786277264, 0.536329600942169, 0.409070388707626, 
    0.249500441689691, -0.0356342370866812, -0.0312283563556586, 
    -0.0252234230511371, 0.110302371794501, -0.135497723886794, 
    0.228921779944464, 0.0582481711215688, -0.0136395273411079, 
    -0.121214477371929, 0.0761414546062776, -0.237429565725894, 
    0.0162273713486294, -0.270621788391599, -0.0942891570638569, 
    -0.153611686916467, -0.140085240532682, -0.0850164770145143, 
    -0.146099002038274, 0.0180432287332299, 0.0673586238436092, 
    0.0754844458556148, 0.0838197777988415, 0.0828012066511241, 
    0.0785881267158755, 0.0715185381653428, 0.0888161523000364, 
    0.0858238888754154, 0.0476624408046648, 0.107218159568093, 
    0.121093827771702, 0.173270153117313, 0.259561436732307, 
    0.204607025716833, 0.0620422535250203, 0.200592157540782, 
    0.403416646364532, 0.149958875960914, 0.133005957536687, 
    -0.245617180718622, 0.445665635800166, 0.328685542946941, 
    0.0939909580542025, 0.406840423165926, 0.382393301263001, 
    0.0397784764765722, -0.419015090920049, 0.11228089871485, 
    0.713464266547905, 0.3765724224716, 0.183759484121689, 
    -0.0752024395045614, 0.687580849383548, 0.216358164955819, 
    0.0939015196926704, 0.130051053697584, 0.198480283669588, 
    0.518844859845251, -0.0293962115907411, -0.109714678557119, 
    0.042659898771571, -0.119321055925697, -0.00556407718309455, 
    -0.255803159778642, -0.0884701222780708, -0.0313862362221835, 
    -0.0987736187762266, 0.0956848736541078, -0.159091089126171, 
    0.183287864578805, -0.108861377961518, 0.262745072556887, 
    0.397668761432092, 0.0766969860596435, 0.0531269856034283, 
    -0.279261358603758, 0.341342883428106, 0.369499985227758, 
    0.124854603677547, 0.0301464595440047, 0.659458865800263, 
    0.162198254239207, -0.240765813597155, -0.0702858284194624, 
    0.903072708671252, 0.0105213039491755, -0.331540623408324, 
    0.191452614041177, 0.623802011962075, 0.0304524675633506, 
    -0.0274659385644192, -0.0808458949411992, 0.0244240855333801, 
    0.37634801050786, 0.496762375711358, 0.198285017978828, 
    0.0177852615472537, 0.0542253358626351, -0.224619109049838, 
    0.224849869920547, 0.537029544036071, -0.000996929740536265, 
    -0.154873284825392, -0.0786464574232778, 0.240347667729769, 
    0.260966973916413, 0.458644610854575, 0.275105582020342, 
    -0.180220744948895, -0.346619635749782, -0.117832384002549, 
    -0.176111669835244, -0.193015410808604, -0.122823089501205, 
    -0.201656820919783, -0.130826142677134, -0.160912175827033, 
    -0.131283971222124, -0.133931564437236, -0.0159136989034647, 
    0.0446531425456175, -0.079296496592966, -5.27624117986625e-05, 
    0.0523748840425638, -0.0409383157086661, 0.0577024553253584, 
    0.0308748428600896, 0.0481870663244468, -0.0544949663408842, 
    0.0267865150934412, 0.0736253634147995, 0.101914926136008, 
    0.137022633760096, 0.107264332120131, 0.0233519759669128, 
    0.223841055086688, 0.189073517882841, -0.00225404663985949, 
    -0.0572977083288017, 0.136573650678983, 0.239445282355364, 
    0.31177324936992, -0.0785154149962983, -0.138835856105857, 
    0.60710540264887, 0.553917197852442, 0.508944078388849, 
    0.393122397081899, -0.0623963962227881,
  0.18567686359238, 0.0852757202952771, 0.0812084289911298, 
    0.0813225584185794, 0.0784357617506422, 0.0727909764428197, 
    0.0890601111536808, 0.106134342784649, 0.101017909718538, 
    -0.081621213957019, 0.417176418664981, 0.141912123575486, 
    0.00847937805447749, -0.117677281520826, 0.477081613796178, 
    0.246770129765624, 0.0638683133879719, -0.0769077626931036, 
    0.217982356943979, 0.24447267303022, 0.478375870390556, 
    0.398126501081958, 0.257456398555859, 0.792689453970009, 
    0.066717809821474, -0.270132686241443, -0.0541184990427965, 
    -0.100076728786091, 0.469169806192731, 0.0581334168009089, 
    -0.0469531807231271, -0.170236048464501, 0.0994679800831135, 
    -0.102816794364475, 0.0498780483773215, -0.177928017417207, 
    0.0289247346238714, -0.137243733052907, -0.00405107928645115, 
    -0.167123003563744, -0.0142962743202632, 0.0423710118179478, 
    0.124692664417136, 0.320008172951929, 0.249472351717819, 
    0.0652865343485971, -0.0978376545307475, 0.468064197322981, 
    0.360293008534981, 0.14202927968513, -0.0992524139295244, 
    0.655958310599292, 0.445523971388971, 0.133329205334994, 
    -0.230762488279871, -0.0392287526484603, 0.595249590659462, 
    0.308590884873154, 0.0179526240668672, 0.536547401050688, 
    0.477632116406626, 0.168967191510518, 0.0215005275629114, 
    0.408960287596661, 0.163030788911651, 0.0363872372029897, 
    -0.00893760314151086, 0.00614062153882991, 0.178658380457281, 
    0.364106620901153, 0.180145713293493, 0.0880267925540426, 
    0.0764730529274358, 0.0247793147463714, -0.01328939210126, 
    0.0356902780084209, -0.090090412489283, 0.044677933511251, 
    -0.0956236021508282, -0.093911406252843, -0.0364226645712481, 
    -0.0178761975637146, 0.109392066347278, -0.131688026893046, 
    0.068867928512952, -0.190842874019179, -0.0451996225342939, 
    -0.110661659026575, -0.0282028597372375, -0.143294290429696, 
    0.0864601369615907, -0.0557105005328717, 0.0938147671750754, 
    0.274107339131463, 0.117435843146104, -0.0186109268858341, 
    0.158831267300739, 0.260255721693722, 0.0913197108198169, 
    -0.476692983428089, 0.361552757809515, 0.546336068815036, 
    0.339432654472708, 0.135159580979349, -0.324108350128526, 
    0.153716950454243, 0.302941860543209, 0.186580524191484, 
    0.806677776448824, 0.601243468740911, 0.389364587553176, 
    0.548985779704566, 0.196314403250997, -0.00898650447855226, 
    0.0690631066077056, -0.193150678052743, 0.0635941963376165, 
    0.0283182082759577, 0.608853683317566, 0.331515104475383, 
    -0.145745070836336, -0.109381888868965, -0.0880841531694517, 
    -0.107906086191129, -0.00578059820742199, -0.0364643531873291, 
    -0.124873578961452, 0.0919648771147504, -0.166587684814483, 
    -0.124921110912484, 0.0119174383166497, -0.129613657446251, 
    0.0322751453059495, -0.0622812573328522, 0.0187650321392222, 
    -0.155761981080211, 0.0184348053171943, -0.0972734680137548, 
    -0.00354399582460618, -0.17023364288301, -0.0512400530434915, 
    0.08403362688526, -0.011836940592039, 0.164932564407835, 
    0.177069994679476, 0.0484909082255771, -0.0455943837686143, 
    0.0727627019946667, -0.0747095485205244, 0.402296413415922, 
    0.40282746139745, -0.159562219118761, -0.0369015578953419, 
    0.491751287787117, 0.548158818066758, 0.324997473332481, 
    -0.236501888685461, 0.416039840647755, 0.462782057996521, 
    -0.0294666002303825, -0.261690564413452, -0.0962898585691191, 
    -0.0579724255622542, -0.176441332537396, -0.0242570119958472, 
    -0.183619644583351, -0.0506523927762861, -0.118773333507726, 
    0.0212396717494076, -0.144785140068891, 0.083141280039214, 
    0.0426858831791401, 0.0748645028293238, 0.0833286839050417, 
    0.0757124674288181, 0.0137524704116912, 0.0583152986846276, 
    0.0290844354112606, 0.0531857656037521, 0.0942447192405143, 
    0.00524478473790056, 0.0790182417820478, 0.209178337252309, 
    0.182119201646586, 0.233427507867113, 0.176462568057488, 
    0.0102653831468143, 0.416867247494159, 0.288613450122264, 
    0.0886993631621214, 0.506669696982033, 0.372756232957996, 
    -0.215985070122256, 0.175044848665144, 0.542877700305111, 
    0.614792901842108, 0.242179173828803, -0.359642808502672, 
    0.1959531340914, 0.583573695426776, -0.021059357941191, 
    0.00939544100783962, -0.211302857681228, 0.214652162215984, 
    0.399741230293694, 0.110086946131934, -0.00470780727042866, 
    -0.0675985635425361, -0.0475334064986463, 0.392695021022401, 
    0.218210738982206, 0.0780067028845949, -0.153585650429483, 
    0.202920969449738, 0.266719390376235, 0.117046443257171, 
    -0.0216076922172802, 0.263320001915618, 0.145616228972852, 
    -0.0175751980375139, 0.0608466321411514, 0.311017566490605, 
    0.183573919718755, 0.138638809178385, 0.0871379758185552, 
    -0.111936437019521, 0.15036267353888, 0.420871953199458, 
    0.00840000057239004, -0.00228030940418665, -0.158969449080529, 
    -0.0364934453283376, -0.0867961754135172, -0.112234124209177, 
    0.11044982493655, -0.121308797444916, 0.0451038567534812, 
    -0.0743018343617114, 0.0397623289906483, -0.154469585570471, 
    0.027881233748519, 0.0825487193705816, 0.0518188519063901, 
    0.17495448111556, 0.280888243319185, 0.135619288226105, 
    -0.0535880094864655, 0.147648095419285, 0.462131874138907, 
    0.1517413449938, -0.205398827299634, 0.255888347422961, 
    0.499941650529552, 0.130047085588116, -0.0389461298910506, 
    0.30974111820251, 0.665754825124665, 0.383664832481591, 
    -0.157548640642533, 0.635780651933143, 0.731317279967925, 
    -0.170380194169774, -0.153956710627673, 0.0841199850754909, 
    -0.0886463983666324, 0.342491022674491, 0.174440575795059, 
    0.0853716140643788, -0.0592998757031997, 0.0285990541075329, 
    -0.479530932028263, 0.063905403994635, -0.341299286755113, 
    -0.383968805925266, 0.368262089820795, -0.405982031720176, 
    0.0904565456589101, -0.512691231828555, -0.202565884790216, 
    -0.155029986288469, -0.0657392289579205, -0.00510195419374322, 
    0.127388670368261, 0.0936099055557852, -0.0351537983532192, 
    0.116752305861343, -0.0232545086937422, 0.016420237771063, 
    0.0640563524570061, -0.0792262479411173, 0.0201314880603257, 
    0.0495498806917655, 0.0678357873322453, 0.0960230971749523, 
    0.10740294683199, 0.0944324282662196, 0.115050376025224, 
    0.121094572331326, 0.0343916358870124, 0.138918136721913, 
    0.362649878920915, 0.149354813390974, -0.173937142753062, 
    0.349028763621844, 0.425405527049314, 0.150910099425524, 
    0.137615318119798, 0.618971679105318, 0.217665755579176, 
    0.0411902793109687, -0.0743882249679658, -0.374778985031949, 
    0.62414588910306, 0.593260611023258, 0.366298914532645, 
    -0.425446345289677, 0.50546109567263, 0.452435624752433, 
    -0.0117171978799833, 0.61986990413389, 0.367556454147801, 
    0.0469545766567565, 0.0453330868063578, -0.175917167947339, 
    0.195049349680392, 0.079646343153182, -0.266469163057104, 
    -0.245521151814257, 0.0347191711292366, 0.241319815467255, 
    -0.195761239881023, -0.0219520103387038, -0.0634985860845625, 
    -0.0630164699498065, -0.0510684878593532, -0.0443402342212635, 
    -0.0683828881834347, 0.0568561638248851, 0.0777841627926079, 
    -0.14347715128668, -0.191376128933391, 0.459113581545659, 
    0.191162523646023, 0.0496101988389328, -0.0974834033760302, 
    0.00532293101913853, 0.0645141060490233, 0.476727225609947, 
    0.554601047993156, 0.0915021436877132, -0.22225189171047, 
    -0.0149480718089047, 0.573528402206467, 0.189592091466538, 
    -0.0836308296525506, 0.317620273145932, 0.348974473348699, 
    -0.00578747023888473, 0.253696036626018, 0.555796604166254,
  0.412360203906566, 0.277916010638962, 0.173892332040818, 0.112668230385335, 
    0.0636523356189254, 0.0295873119646686, 0.193071954514709, 
    0.425895998675875, 0.120906154342581, -0.22447840624594, 
    0.0648177094614105, 0.226355699356622, 0.388419401404344, 
    0.622997046285264, 0.27113943375366, 0.101945736640013, 
    0.290313346821353, -0.569756406746062, 0.307730283712868, 
    0.715391204273173, -0.0825637500183287, -0.00931883053607188, 
    -0.306022733760128, -0.119159024676914, 0.729776020767871, 
    -0.223820178320419, -0.376510908349516, 0.106892609321554, 
    0.577872591164567, -0.17076502780933, -0.054993660508589, 
    -0.227228432581564, -0.0925431042765395, -0.0943897607155339, 
    -0.194495406674335, -0.0799140770130897, -0.167126073074541, 
    -0.0993262410266329, -0.0596204246109097, -0.0976469401935853, 
    0.00627179337081089, 0.0369481222576078, 0.216960685853284, 
    0.165847930535565, 0.0743200188065429, 0.115893262304375, 
    0.212196430692865, 0.165801477853171, 0.0871364575919608, 
    -0.00879328858460977, 0.228700863634909, 0.212962339176977, 
    0.0604618137598107, 0.15847823622879, 0.334808814822001, 
    0.17623634423556, 0.0443087020855561, 0.234734430336254, 
    0.28999946321204, 0.109039388772918, -0.00304295219701742, 
    0.0245605549949972, 0.0451563129923873, 0.0231556092176145, 
    0.0640407268089794, 0.021394181305515, 0.0338933614185798, 
    0.0533913635206815, 0.0542220414603379, -0.00929205628031474, 
    0.0561722054560565, 0.107942275260653, 0.145116911735709, 
    0.147646814384171, 0.119455198892574, 0.184019781557857, 
    0.309120517591123, 0.169007203659957, -0.0179880886363055, 
    0.0501231824980979, 0.453118595226096, 0.195684358387809, 
    -0.0500432049152647, 0.490993542105814, 0.51968616165586, 
    0.190087856381731, -0.0965244611107588, 0.289590897305712, 
    0.343830693189173, 0.116004383659587, 0.444549791196083, 
    0.382634671230891, -0.0275266107490119, 0.0963868180117742, 
    0.551981854603006, 0.130449258764203, -0.0216217913138306, 
    0.28175773503113, 0.3091410728107, 0.128760513455268, 
    -0.0524388396980728, 0.0521378522137652, -0.454610622350669, 
    -0.0663777229963009, -0.0864940631737538, -0.299413793074489, 
    0.153325052048685, -0.0971195659603943, 0.141786914353366, 
    -0.192764233212238, 0.106446245066981, 0.0815576678786445, 
    0.0792320126974657, 0.104257338644264, 0.111138372561644, 
    0.066290686920327, 0.0952401340175642, 0.128345843553897, 
    0.1002651312098, 0.0287261294800896, 0.0796237322979458, 
    0.109537827862924, 0.152806230978168, 0.180188000372693, 
    0.123139841808674, 0.120224732722903, 0.300454670427645, 
    0.227584967240643, 0.105454443600633, -0.0605797930942832, 
    0.578510486323163, 0.0827773484745468, -0.140280648240425, 
    -0.22672174495094, 0.590890981939032, 0.444233163275091, 
    0.0809766401641578, -0.0979559456270457, -0.124295601475772, 
    0.565623293668469, 0.169263266706394, -0.058904872045321, 
    -0.0919266594019654, 0.460921868137249, 0.44991142112804, 
    0.0766481750142114, -0.328984594774317, 0.280344171724707, 
    0.341880459165671, -0.382774854523461, -0.199768013395665, 
    -0.0789396689693083, -0.170551942684739, -0.0780690725579444, 
    -0.155594529690745, -0.0335158035831514, -0.137515529903419, 
    -0.0463270999529188, -0.0866013696781164, -0.147335699169244, 
    0.0668805814734759, -0.0830385351457717, 0.0511360590721584, 
    -0.0585461809693306, 0.0106907594784152, -0.0131627744756369, 
    0.0613068215720883, -0.0359961946303872, 0.0752477665232528, 
    -0.0549122765041333, 0.306250160146266, 0.120825023821259, 
    -0.0395835510277516, 0.0292851996814643, 0.239769624031053, 
    0.24246828058634, 0.299349064398824, 0.306707014323317, 
    -0.00713446548803015, -0.248395758810802, -0.226087092643747, 
    0.788747375011168, -0.00529891402645841, -0.18962702834168, 
    -0.0391684791869804, -0.0733438400681344, 0.290465486329608, 
    0.977780621063489, 0.443856142851292, 0.0181855381313953, 
    0.616594067359754, 0.543679535308239, 0.191398796435057, 
    0.290225940734227, 0.264512386947983, -0.195489807631848, 
    0.104511367562859, 0.188333184621262, 0.377435385613416, 
    0.514156000052313, 0.0971359595205102, -0.0383768782804454, 
    -0.0394259743843152, -0.126291314483189, -0.041900992133368, 
    -0.167529459051378, 0.144547362996587, 0.208588434435773, 
    -0.175647429916678, -0.169882377922923, -0.0811383044954655, 
    -0.189141114780923, -0.126106039707182, -0.0957488400951366, 
    -0.214669247503095, -0.0809098953384299, -0.12434619760642, 
    -0.178753069993264, -0.0569798863789699, -0.208841416377607, 
    -0.098876653239978, -0.0925593432187443, -0.0314064227501151, 
    0.0906137981379417, -0.199361945439868, 0.0758111108949163, 
    -0.162410832949046, -0.0870451695224366, 0.00311361547540118, 
    -0.266486011575912, -0.0373278050022148, 0.0388373954135722, 
    0.0484034606352577, 0.0636818587143669, 0.101238218435426, 
    0.0773196210375702, 0.0580112042494611, 0.136094169995555, 
    0.124165187553806, 0.199034496864649, 0.279914458963112, 
    0.0198182137851442, 0.253588425161942, 0.448934153594343, 
    -0.0730248861245152, 0.46745790085444, 0.772722641791093, 
    -0.259658486990381, -0.384019200343337, -0.126760875098599, 
    0.569282465541189, 0.355735572326686, 0.356786899547025, 
    -0.0683218946845297, 0.662908106889334, 0.156990359749671, 
    -0.0412975740526403, -0.162860924481978, 0.601103262478266, 
    0.372485775347361, 0.149188562482895, 0.159728693709976, 
    -0.084912845721436, 0.499054726335962, 0.207460403567808, 
    0.206203232227406, 0.204190074328776, -0.231978522297059, 
    0.139649029278148, 0.535506690144441, -0.100770427425442, 
    -0.00806113515480972, -0.166658993566183, 0.0139097493497654, 
    0.0603944674865805, -0.0443259159593599, -0.135364877580777, 
    0.0266694923165688, 0.0757692816592302, -0.0803487745570841, 
    -0.0251492345810078, -0.150718849728499, 0.0924208415371278, 
    0.0578359123504012, 0.197433744326775, -0.258419333933345, 
    0.189478139889204, -0.308463459474707, 0.0110879073661711, 
    -0.232926089661374, -0.0547937217779351, 0.0124659429005699, 
    0.00929540793447185, 0.0150473997612931, 0.0326630529230769, 
    0.0237327546828275, 0.0117412046399443, 0.0343398994885858, 
    0.11681561873623, 0.0511743400226158, 0.614450207154468, 
    -0.0767992508087655, 0.0342950464384804, -0.306890770634068, 
    0.244815782350675, 0.385044910901003, 0.367225814539725, 
    0.553738350789994, 0.322802434921153, 0.0327983395334465, 
    0.162538480057021, 0.422321812588843, 0.167414393767696, 
    0.0867776285265783, 0.0988045335816638, 0.017938939104394, 
    0.00684356025212435, 0.217580820549415, 0.0360765684722953, 
    -0.019058347005343, -0.02347680276102, -0.193807478471969, 
    0.10113943789864, -0.0949457264192421, 0.076575977774625, 
    -0.231839053060477, 0.0293753659492233, -0.0727680111548263, 
    0.0911275844675357, -0.317901628776698, 0.0517938301107556, 
    -0.205078554186256, -0.111542983787317, -0.149138061819447, 
    -0.120864367535608, -0.149670437984236, -0.106925215443937, 
    -0.102968316874675, 0.154985382979209, -0.466945806311406, 
    0.3729485172294, 0.407724698002013, -0.130908114954738, 
    0.112328920906358, 0.0628565907228197, 0.12658772983017, 
    1.01305850778409, 0.4899810281893, 0.115047183061652, 0.0740128167817391, 
    -0.0879127004034378, -0.0972665875042669, 0.051833321574049, 
    0.277336786767269, 0.508150259098175, 0.566692534099008, 
    0.399161458505923, 0.216568306117291, 0.216286057211275, 0.448947040784792,
  0.0744726473094795, 0.201146339147381, 0.132160806051256, 
    0.00382093262210348, 0.320345600065234, 0.239775743067049, 
    0.151185001583568, 0.469311200889731, 0.288416854043644, 
    0.015574179041653, -0.0710863743283663, 0.0120822652260755, 
    -0.257349118080628, -0.0428673405075296, -0.101056220797633, 
    -0.169639374590542, -0.0222504696293133, -0.0076698069245581, 
    0.0683704782149634, -0.210489553495655, 0.195823905763364, 
    -0.0308359300749556, 0.535704009200864, 0.243962940087418, 
    0.100103444908268, 0.130695301836589, -0.308945938399044, 
    0.222107355927352, 0.424713907338859, 0.199795430805495, 
    0.116776534208861, 0.320282180114694, -0.033117609669913, 
    -0.0725863273048958, 0.812994645037703, 0.311092657338628, 
    0.107460782871325, 0.970722918331459, 0.323393075310911, 
    -0.00229454709726511, -0.117513498963701, -0.208352628636099, 
    0.0895027180811631, -0.114382350294785, 0.0871838092948366, 
    -0.118090900413888, 0.1043728736257, -0.130206910101175, 
    0.120119136301853, -0.154603649637325, 0.143427673176706, 
    0.00836851201535062, 0.225249542021905, 0.261215018823611, 
    0.090364867133225, -0.0702737425624521, 0.285737784739916, 
    0.232666126494184, 0.023584461569677, -0.26259613135547, 
    0.376833917685584, 0.652576795277947, 0.36748565700595, 
    -0.205114524810279, 0.91081912978117, 0.704651126698655, 
    -0.00866228305312682, -0.0512591298073741, 1.42187292891778, 
    0.191915321155231, -0.0623633035384038, -0.00157828529356416, 
    -0.127243881287814, -0.0626393631141183, -0.0398657698311134, 
    -0.21046413136733, 0.0290639759582982, 0.0448845480137957, 
    -0.250274133608956, -0.0234849696893859, -0.0944843943682833, 
    0.00550651226588612, -0.0885711619821814, -0.0367484042625645, 
    -0.0550953243327739, -0.0459558821330585, -0.0149467007062692, 
    -0.0500236267358549, 0.0461179219360897, 0.0510176709969206, 
    0.3717038787202, -0.00759231691580693, 0.227802601680681, 
    0.527616658304114, 0.0452822887187057, -0.151464277082578, 
    0.148555991687702, 0.346607309538414, 0.0587388625128106, 
    0.0784244315394389, 0.320232761670796, 0.264265071167354, 
    0.190747943048597, -0.162582802811225, -0.0830510651836233, 
    0.64108719508847, 0.232473640406745, -0.0703330520819284, 
    0.835116243887506, 0.281566383957373, -0.070806185778915, 
    -0.0259431504880502, -0.187633441674235, -0.0468109207252881, 
    -0.266301629760756, -0.197453925862588, 0.071116409555721, 
    -0.0851337526522669, 0.117009954949945, -0.211569319678584, 
    0.0164870527805828, 0.109622020309603, 0.205086257510858, 
    0.215715866153587, 0.130979648651494, 0.129945460975487, 
    0.371706699135215, 0.425377242016903, 0.265728866640633, 
    0.154904401131815, 0.22557178499011, 0.382973641774713, 
    0.410130556245437, 0.332762689947281, 0.318747228008409, 
    0.441609062509886, 0.426376925363887, 0.231864386244239, 
    0.198252030385709, 0.549878008097735, 0.354847029193132, 
    0.0426253232232164, 0.320542457860299, 0.544212822182186, 
    0.0692776670767802, 0.0227171604618215, -0.237368450078867, 
    0.438686523385166, 0.344166887398846, 0.0191234917164428, 
    -0.089820322607687, -0.257951403179892, 0.319996119598004, 
    0.37844195914528, 0.0793684058517994, -0.113310867533179, 
    0.0352710499268731, -0.0923215259918496, 0.281235740962889, 
    0.544132855903546, 0.121114955634126, 0.00977898591611853, 
    -0.0169578333324725, -0.0657943071336243, -0.086112480680246, 
    -0.125826188747476, -0.0415067376770845, -0.150330265751158, 
    -0.0584385902312073, -0.127015282342331, 0.0637975428122246, 
    -0.0279024752397136, 0.057597578904132, -0.0105977218835515, 
    0.0422361903823626, -0.0255409051293538, 0.0136199390455976, 
    0.0476357120071538, 0.0987358274988143, -0.0719179656760035, 
    0.0320284587701071, 0.219004182006835, 0.186915658826441, 
    0.0875320671477584, 0.0291965799149414, -0.12885757894909, 
    0.178046726016744, 0.366830801795168, 0.18276884120156, 
    -0.0867437275849968, -0.0474094597012075, 0.638544589269382, 
    0.926864692392867, 0.265560444984519, -1.02006427175169, 
    0.46785485725139, 1.04230872399252, 0.388909770061371, 0.305363997116924, 
    0.521388016865433, 0.0284563792274682, -0.0625302972209524, 
    -0.0590149996753555, -0.140561068303664, 0.0248070663506833, 
    -0.253138094495719, -0.20496969242744, -0.328904253510129, 
    -0.110220625516703, -0.337479250057109, -0.00342034158848273, 
    -0.13706754960389, 0.0573922989408873, -0.175366750930775, 
    -0.0295584559594524, 0.175812212732368, 0.153824042081819, 
    -0.141784623571043, 0.168595005239553, -0.209558459821148, 
    -0.045107498266248, 0.0235114450532458, 0.00813221514521011, 
    0.00050725141381433, 0.0280298553090174, 0.02280721686757, 
    -4.2664576004825e-05, 0.0532209429466629, 0.0198562002856193, 
    0.00104558005050033, 0.143781723243388, -0.101195580161556, 
    0.326031834461525, 0.330523364910603, 0.121239837429078, 
    -0.144817800270395, 0.238055994773678, 0.398992797951516, 
    0.100576215503182, 0.00421347407383886, -0.129876490693392, 
    0.457676473594757, 0.323481505296551, 0.19968106786184, 
    -0.168351240709711, 0.426232697822808, 0.254451415813913, 
    -0.0285974870791802, 0.146667350412908, 0.451184738038745, 
    0.175151209519567, 0.0907042693189245, 0.0845766400812549, 
    0.0838846526893662, 0.0647470863157995, 0.0754785854842261, 
    0.0652804368518938, 0.0595487134316178, 0.0637454625715186, 
    0.111246985498654, 0.162393878085412, -0.0326216831704579, 
    0.148056444039851, 0.362782873387074, 0.305936249376135, 
    0.175190309307366, -0.169561083904417, 0.368304961549667, 
    0.393204569781595, 0.124212775014368, 0.151303288120868, 
    0.326361929722114, -0.127409977556296, -0.259913063004407, 
    0.979275653577363, 0.326508844795853, 0.126763087034446, 
    -0.294879054967336, 0.266400485566619, 0.511830107022557, 
    -0.320349051733332, -0.0338661265838193, -0.136068078013705, 
    -0.0404430397519733, -0.281576126187213, -0.112842572925711, 
    -0.0468520956446725, -0.284589426038014, 0.0837584320193549, 
    -0.11382720853698, 0.10948144242703, -0.0462510607407558, 
    0.0922166705198058, 0.00390777721422818, 0.0682082485826543, 
    -0.0521763139893616, 0.0446763784437832, -0.0152638767615561, 
    0.0406298862817738, -0.205784947523779, -0.00310651725462639, 
    0.000832445359803452, -0.0024653330463997, 0.0806451084707299, 
    0.048134893966089, -0.0237874025331597, 0.016272472503253, 
    0.15760834580553, 0.12063277465161, -0.100437695425633, 
    0.498025453182934, 0.040176182272692, -0.0138752216865725, 
    -0.259409234010019, 0.019698548239425, 0.45241164508223, 
    0.497124389405195, 0.297426890959622, 0.109491292619021, 
    -0.0596704738236875, 0.112066146445415, 0.323618308899052, 
    0.177404279703011, 0.0960672125073566, 0.0788181500639701, 
    0.0748733748832455, 0.070164502322567, 0.0715420934833362, 
    0.0712999009038517, 0.0623426097833827, 0.0557891269446221, 
    0.0695933078869145, 0.0831625595158775, 0.0831768475282716, 
    0.0660134646280418, 0.0695216545653854, 0.0643202454515904, 
    0.0753866967300622, 0.0792927906227193, 0.0709391922469951, 
    0.118444787110966, 0.111759874672521, 0.0970613444856531, 
    0.0938356806947891, 0.175664473880677, 0.152319177551502, 
    -0.0318491833553091, 0.347386941530336, 0.204768986133716, 
    -0.232126276786277, 0.232724438407713, 0.460293627471961, 
    -0.0569310029312472, -0.273826381483675, -0.147040138194265, 
    0.504268495486913, 0.221001288856745, 0.158283766204687, 
    0.747501250643362, 0.368524831462589,
  0.602065443355149, 0.49729671128508, 0.193645981070379, 
    -0.0621333645653937, 0.327559665377326, 0.0614693821773599, 
    0.247137762645781, 0.948280129644939, 0.081072314526915, 
    -0.0990085636772602, -0.188633097491743, -0.227743898646073, 
    -0.0197214668655303, -0.323345499287791, -0.107506617523678, 
    -0.213100790442437, -0.203146845088141, -0.147852317250581, 
    -0.140802662327374, -0.168029064829767, 0.00351981618160888, 
    0.0563614993683837, 0.0260628065119536, 0.0718373306774241, 
    0.136657748331773, 0.0207609364675359, 0.0609134817883422, 
    0.0837564409837499, 0.0785387108804023, 0.0177938714808166, 
    0.0557815732130609, 0.0829419482797693, 0.100971874485626, 
    0.142410298867677, 0.154655853366638, 0.096244139359666, 
    0.0994386983927338, 0.249735306819408, 0.103575689064065, 
    -0.0241512888316888, -0.0614404427595925, 0.334661747989139, 
    0.238330527070972, 0.229075610228418, 0.362027676219361, 
    0.0536044228834388, 0.0512084460993486, 0.686933364051402, 
    0.462858433914999, 0.10541671778674, -0.223534363514655, 
    -0.00884588713011636, 0.432500674943679, 0.276681172281126, 
    0.0996802601834222, 0.0491454219320607, -0.272019490799207, 
    0.319479706534959, 0.380846620689204, -0.324408222113427, 
    -0.235870737585085, -0.217597434565675, -0.0236279393520651, 
    -0.203349153903699, 0.000666597254732448, -0.218369540334506, 
    0.00304816716140299, -0.19117169688314, 0.0384970054941814, 
    -0.174505039850976, 0.103890992721874, -0.0250417749347131, 
    0.0576211549520975, 0.0194844365200303, 0.0648170102478378, 
    -0.0452232343104191, 0.0367934728607133, 0.0204045551111355, 
    0.0404105082996481, -0.0890604598767951, -0.00703188145757089, 
    0.11784152133919, 0.0940372006228122, 0.0641688317008991, 
    0.2253819543266, 0.16710605182297, 0.01767446473073, 0.0410003284284791, 
    0.424289526339326, 0.0468243091191877, -0.11504783394937, 
    0.0322780602393051, 0.536619683001686, 0.166719134615635, 
    0.0598244831791391, -0.210408474413358, -0.169147697803653, 
    0.686950449650297, 0.173827813562243, -0.127491754825068, 
    0.0639913438094305, 0.552009100548929, 0.104401588271161, 
    -0.255280130834443, 0.285453008157506, 0.282230437418854, 
    0.0688406064631481, 0.443429776706683, 0.13642312433844, 
    -0.104199970345221, -0.181496372696019, 0.0404573489998404, 
    -0.156160426941601, 0.0456170151699777, -0.120950793027914, 
    0.0781751172726598, -0.309492586232469, -0.0108162909657696, 
    -0.211295131081061, -0.192528968511579, 0.0156996421660103, 
    0.0749796241795827, 0.099001180615619, 0.182467539705395, 
    0.246237366154705, 0.212090408187748, 0.217308405317846, 
    0.225588898132698, 0.0907733599086945, 0.172338613070557, 
    0.62511452737396, 0.324043529146433, 0.048131299651803, 
    -0.0777366180169129, 0.670778191493697, 0.377108074731993, 
    0.0751846275523897, 0.0224198341703904, 0.7956760966399, 
    0.0951165230997474, -0.243287068327467, 0.113513601724468, 
    0.534758522747508, 0.162189286137368, 0.448012432648448, 
    0.323384287082183, -0.355734211052926, 0.0683974447942798, 
    0.521385323288509, -0.0934493887052994, -0.294108318050551, 
    0.0442600879867486, 0.104158467892833, -0.0494624197043849, 
    -0.0139726252337651, 0.0316991013716366, 0.0751695920439689, 
    -0.219657096966448, -0.134066634153182, 0.0817608123132648, 
    -0.409501835368125, -0.0683883827846851, -0.121637351358132, 
    -0.241450933081807, 0.15015931477597, -0.233776165618754, 
    0.0235025592022306, -0.0207018650070531, 0.121646071030749, 
    -0.205660142942619, 0.0565870829201531, 0.0562825777158855, 
    0.0651305001605949, 0.0715697891078833, 0.0894848848501851, 
    0.0642165025908046, 0.0657891860328422, 0.102906629991888, 
    0.0912208499931537, 0.0325637215144928, 0.0943530453238403, 
    0.123880799624041, 0.135851159867742, 0.17516709375574, 
    0.191784203859258, 0.158809244135774, 0.183171473502821, 
    0.23364785563775, 0.137421867481712, 0.047803569039448, 
    0.403978614053653, 0.269217711155133, 0.0346491559677364, 
    -0.0562643652626187, 0.491878134078557, 0.327642516463197, 
    0.0760758135451112, -0.0858815747748177, -0.0902368342900974, 
    0.516329902294011, 0.382040726946074, 0.188215837356045, 
    -0.223553812959685, 0.371310525973376, 0.458462322702528, 
    0.251196856541457, -0.0297454905643831, 0.644133647314217, 
    0.0561764099981907, -0.178452462649687, -0.11302787008348, 
    -0.275957958854224, -0.0966818546586218, -0.0963375737111913, 
    -0.0676380948614297, 0.0471971415287899, 0.158639037080191, 
    -0.249729760208864, 0.223238066414515, -0.221994834022915, 
    0.0942896750949881, 0.102573362577359, 0.014541524714849, 
    0.223157806410794, 0.453637166384925, 0.231518067309869, 
    0.0248724413610363, 0.0950836699163158, 0.445565030794281, 
    0.211839344836573, 0.0920980015421751, 0.139223354636048, 
    0.0770320747038595, 0.0919725859225575, 0.106494495933629, 
    0.0769465130990746, 0.0746852415818736, 0.128356515955303, 
    0.255099210999664, 0.151821041555942, -0.135404230416232, 
    0.31369296397461, 0.33904434757966, 0.113222610935254, 
    -0.145000679118237, 0.199615577097984, 0.356356253365316, 
    0.229067440001366, 0.221359860599949, 0.20089126818972, 
    0.430431987069014, 0.422195874285385, -0.156906348154196, 
    -0.460564064085149, 0.4389024492684, 0.871058703575996, 
    0.433236589519058, -0.0217850967687771, 0.642277902922907, 
    0.367138415375572, 0.0516389869253806, 0.0540473908635485, 
    0.0243364343546792, 0.0219115071625864, 0.0639405023997336, 
    0.0198194118102499, 0.00745541887175, 0.0161518613568231, 
    0.122298664360241, 0.0928640414746128, 0.104653315329171, 
    -0.124893335743026, 0.307271057949538, 0.344351715745672, 
    0.140763735983751, -0.00861659053857655, 0.150604658474459, 
    0.137001498689184, 0.0662868008909435, 0.692439725752431, 
    0.322219226487329, -0.0165017414390661, -0.0270528019231673, 
    -0.1969760824455, 0.110186862027366, 0.399244161053235, 
    0.961207427578014, 0.318274044693567, -0.185751566651751, 
    -0.0816654944100267, -0.0772201290177887, -0.231106637703385, 
    0.00383211066956907, -0.227034113194881, 0.0723444573663448, 
    -0.205280577732864, 0.0921421269111316, -0.201528420119645, 
    0.0672107148885999, -0.216702220584763, -0.0144439959218871, 
    0.0974169299352104, 0.113888736868565, 0.169303938654015, 
    0.248324363237154, 0.163037811704797, 0.0745591948386295, 
    0.261638435944508, 0.230551230068906, 0.0564104723801839, 
    0.12910706016564, 0.344206727548043, 0.322982872406966, 
    0.219746204905734, -0.0438926975907869, 0.186917286223751, 
    0.922450461623284, 0.153320161383002, -0.110072892471241, 
    -0.0700632207298098, 0.487899327773376, 0.361848359584293, 
    0.279372904370039, 0.105802569033159, -0.0729435944353814, 
    -0.285944584806413, 0.174173049574566, 0.595353255514353, 
    -0.0888903004198811, -0.0222475616531241, -0.284967490966299, 
    0.124886217049832, -0.322443565170895, -0.10975354103956, 
    -0.145948117308064, -0.17851040660712, -0.0194113858825642, 
    -0.150275894279789, 0.0724953439109264, -0.205137517212565, 
    0.0250484398204081, 0.0896684012977325, 0.105286778358877, 
    0.142347446047779, 0.158573938499045, 0.106673137250816, 
    0.0853561224749978, 0.191464858946334, 0.156756430294302, 
    0.0476884396032854, 0.0163680830412366, 0.217704986599363, 
    0.283485143635513, 0.245568620718199, 0.212085291691836, 
    0.169342789295327, 0.423397227048976, 0.356287512040984, 
    0.0457398867340953, -0.0547253281491278,
  -0.0935112927891758, 0.0213576451439944, -0.00393436998229388, 
    -0.24547359005166, -0.0562437169542829, -0.0232080659239305, 
    -0.0367839679840805, 0.220968505197637, -0.19160044751363, 
    0.0320161505770967, -0.104334984645621, -0.0294379538919421, 
    -0.0700205843842343, -0.0488021496136752, -0.0776479276089132, 
    -0.0455193813951817, -0.0550427103363985, -0.00544073533016701, 
    0.165375527214295, -0.189282211235749, 0.0764397061436906, 
    0.307706002296182, 0.22540493666774, 0.0418645986697839, 
    -0.059064670291917, -0.223094822756725, 0.394094476481544, 
    0.30930469124844, 0.0860196235865492, -0.244249830155301, 
    -0.164842870449866, 0.247679152355887, 0.740246709594599, 
    0.371710925138489, -0.201723743085016, 0.359490116600897, 
    0.707463627670329, 0.225976170643289, -0.0976859337175009, 
    0.0945658603297052, 0.587406198492392, 0.200200632149235, 
    0.0203267179899892, -0.108452122104007, 0.34594967021768, 
    0.342495761305583, 0.087810907664647, 0.0103733643542828, 
    -0.122342173991292, 0.373808424406211, 0.193255238297927, 
    0.0696995901801925, 0.261032134513432, 0.213454889572266, 
    -0.197361770415926, 0.141944813559083, 0.380152085785752, 
    -0.0205335922747255, -0.145735168299504, 0.0698643629066569, 
    0.217218033004397, 0.0163934234641397, 0.241002720965098, 
    0.233979303019183, -0.156348204387269, -0.0820935534182708, 
    -0.0664610009808588, 0.236889753269743, 0.0575894373314834, 
    0.0358268723676117, -0.168802271509591, 0.0417524787641531, 
    -0.184956989511685, -0.0274555441280983, -0.141373137900173, 
    -0.105420761327514, 0.00699215939840343, -0.0874562859619397, 
    0.0614323230123117, -0.14444623585078, 0.00272126636383824, 
    0.0633481927947656, 0.0848885187227332, 0.104839001607594, 
    0.113201523979056, 0.137177901333759, 0.193652812937469, 
    0.0989365398957895, -0.0854675001220713, 0.0297295327965228, 
    0.464420663420085, 0.112528796741596, -0.187018288180178, 
    0.472016976235511, 0.559470606423006, 0.226772596864243, 
    -0.0506333286831929, 0.491715462910815, 0.413314059057619, 
    0.467372984336142, 0.357296718200388, -0.223090743688864, 
    0.454802505603317, 0.39563085676394, 0.0632160511412328, 
    -0.16836450379941, 0.582014387595994, 0.373258636789914, 
    0.118495609741042, 0.387126603509635, 0.373740168768572, 
    0.158778692775584, 0.0723604642728356, 0.0657714212634521, 
    0.100242371464422, 0.0792743114341167, 0.0434886223519931, 
    0.0965712099459624, 0.0768161374964472, 0.0934577396437913, 
    0.205848261740837, -0.166181363429464, 0.265134411344292, 
    0.372580864952988, 0.380771420980692, 0.230000790671337, 
    -0.228423822144024, 0.0307484788442227, 0.690900473130339, 
    0.168204129231174, -0.334879409274023, 0.594697265196046, 
    0.413143188297012, -0.305108685528475, -0.0822633651857823, 
    0.962293308572741, 0.047435688353457, 0.0410316349759347, 
    0.404814720624268, -0.443536839954104, -0.501716995288648, 
    -0.181378465981062, -0.192688506473958, -0.374684782389353, 
    -0.0709494924972333, -0.313114327977767, -0.0418149316266767, 
    -0.145247630631689, 0.201148374130824, -0.378529997403059, 
    0.00798161214238091, 0.148806593899708, 0.193461867319565, 
    0.137693143366125, 0.152618901872715, 0.158516368530521, 
    0.19538570232425, 0.170853059057193, 0.1806853164294, 0.0716677786287424, 
    0.0538151066819517, 0.0682767196309874, 0.0538832738928796, 
    0.0614376168828975, 0.0626691052100367, 0.0561667899284591, 
    0.0580862595633207, 0.0899804646206356, 0.106318580872398, 
    -0.00446878048374394, 0.178651271298516, 0.190746158871593, 
    0.0388022464289652, 0.0159156268587483, 0.371259902782388, 
    0.229329845632077, 0.0700833152270254, -0.0818885457240925, 
    0.2238764295201, 0.325817711165111, 0.185193762728366, 0.133167530118472, 
    0.130918847862402, 0.132941951847439, 0.134036089102193, 
    0.130611501171144, 0.153859296065419, 0.188606951837324, 
    0.140159062192045, 0.0476068085141164, 0.207606872244875, 
    0.295373912295793, 0.141639813131673, -0.03002177151953, 
    0.172873644820309, 0.369007624331553, 0.247228474573994, 
    0.187940947669425, 0.178999588267986, -0.273680787740057, 
    0.32677991515215, 0.460405231176839, 0.37051244005933, 0.224580557943055, 
    -0.0196571305241628, 0.29484965690105, -0.0923772389161333, 
    0.263557828393462, 0.944331145449943, 0.126161078033329, 
    -0.109797684081911, -0.0607545523891601, -0.0140653926112713, 
    -0.0266927817089961, 0.0101721192242086, 0.143449921300107, 
    -0.126609395173315, -0.0676709053519623, -0.125378371010795, 
    -0.0309355060461361, -0.208534719503285, -0.11941945445347, 
    0.00869900192979266, -0.134950754776154, 0.0862719483544141, 
    -0.111177345482104, 0.0691046780119814, -0.0927605186390602, 
    0.0409661949702185, -0.153582128843522, -0.0357012927122011, 
    0.0781652878361712, 0.0633768364638966, 0.0564689211541997, 
    0.181390153041856, 0.108134458037323, 0.111339904942527, 
    0.375041210142727, -0.0349170711244824, 0.0333610031551894, 
    -0.371522166295151, 0.178281886937017, 0.536218771858418, 
    0.296194354425968, 0.0421423763926759, -0.166393542277074, 
    -0.292521011598676, 0.423582154069509, 0.465150136587362, 
    0.345850608604397, 0.278974275795265, 0.108966539328204, 
    -0.0511999769331525, 0.508427128594865, 0.317222255377088, 
    0.0623128483629465, -0.0829957682860495, 0.109864636800933, 
    0.332593229121849, -0.0205346981413508, -0.0573834574755957, 
    -0.140916971639434, 0.0616478886890744, -0.0914190290044647, 
    0.0634585955902717, -0.122852244548302, 0.0704124871338893, 
    -0.062774069517702, 0.152831938365751, -0.122509446648006, 
    0.297070238471604, 0.13272695037854, -0.0763011607756877, 
    0.00594082170291259, 0.440197443869301, 0.140781876581212, 
    -0.0511811911206588, 0.197640941900422, 0.283751249357904, 
    -0.129063775043991, 0.253518884610797, 0.623978712823652, 
    1.00239476222915, 0.255409904851107, -0.33876929655107, 
    0.0281222013770304, 0.525629376033132, 0.0742680630619164, 
    0.761677094085251, 0.689956863105066, -0.0198166559517179, 
    -0.0405053321866979, -0.115237533893499, -0.0799154167363479, 
    0.0869839428183277, 0.0846837380082206, 0.0351342960800618, 
    -0.137311868301098, -0.172614783293823, 0.118588353855302, 
    -0.228580886556873, -0.0302256444671315, -0.101249926844715, 
    -0.138008719391621, 0.0405255394399304, -0.142992094432959, 
    0.0243627391397459, -0.0566877615769937, 0.0863887903038305, 
    -0.127541182029243, 0.0460619171519884, -0.00708794712311651, 
    0.0145148355865158, 0.00237704950816237, 0.00514091009178215, 
    -0.0270854304157441, -0.0395449654720024, 0.0383448226885553, 
    0.0566040647727994, -0.0157666491176443, 0.197249382011408, 
    -0.13514771069527, 0.24239870318505, 0.376972046285911, 
    0.150289986915869, -0.0434709305067515, 0.16715842439658, 
    0.507479169331392, 0.052687511900385, 0.350517379408603, 
    0.53197635354168, -0.343137511716988, 0.234341446345574, 
    0.606887460391703, 0.362764371555865, -0.468987994262149, 
    0.794546307771488, 1.02817792375636, -0.0159969154138196, 
    -0.0414488808924864, -0.230965907923835, -0.067064543533618, 
    -0.154823930534648, 0.0303127201822067, -0.225019980073385, 
    -0.0206408091187226, -0.165705544841426, -0.00566545519461129, 
    -0.316830748401995, -0.220310691425773, -0.110389229135029, 
    -0.0973131128542001, -0.0904569849454426, -0.0385836843399538, 
    -0.08113269216242, 0.0345928449928948, -0.0814808618842545, 
    0.00918660533090412, -0.24317006271406, 0.00408847158672992,
  -0.140336405141983, -0.16105561308686, -0.0759167445356112, 
    -0.131816059768582, -0.0148466635017996, -0.14934403348621, 
    -0.0114727634095062, -0.153095714016681, -0.0875100916178968, 
    -0.135392277323138, -0.00661742362250972, -0.117843441512224, 
    0.0619024748223226, -0.049019096382363, 0.0817952200790488, 
    -0.138492402089887, 0.0587253852494484, -0.106123020430762, 
    0.0280326698307991, -0.191190304622827, -0.0454747812141964, 
    0.0620042042215363, 0.0654212243764068, 0.0760433499688061, 
    0.139560233726123, 0.0986852585982301, 0.0449463331214257, 
    0.207802249537899, 0.300363726590723, 0.0861424791003179, 
    -0.211943528774651, 0.0745211115250677, 0.594181219198661, 
    -0.0205143156545641, -0.168252650498027, -0.103499878704876, 
    0.596934612893604, 0.160685709782208, 0.0599091590406558, 
    -0.135695320377346, 0.0278347480351182, 0.427820542864945, 
    0.37659652285371, 0.094948497298356, -0.0242456833300476, 
    0.0995981971626205, -0.329878006911699, 0.0926586115353449, 
    0.521356231464518, 0.169178893017627, -0.106084063200872, 
    -0.133166820189462, -0.231506907617607, -0.176628866394678, 
    -0.0979163941948642, -0.199455013588938, -0.031261226537854, 
    -0.180160577388008, -0.000203280352423146, -0.132228632178296, 
    0.0877564143554115, -0.161959833108489, 0.078733335013585, 
    -0.130530227366582, 0.00127349019638273, -0.0897109859566596, 
    0.0193991183432187, 0.0436460180036583, 0.112140585326284, 
    -0.221429374079286, 0.0619310809566004, -0.040048486267127, 
    0.0531841061482435, 0.0113854341575661, -0.0215851803103103, 
    -0.0979735164324211, -0.00912161356194022, 0.0934632581034942, 
    -0.081072034191875, -0.489550312960167, -0.198154839879716, 
    0.682814217665447, 0.0385754597652237, -0.013554101403336, 
    -0.144879823063615, 0.118126898296065, -0.180228107795131, 
    0.536947068411759, 0.783690028607066, 0.336221982945439, 
    0.126328305104103, 0.167515378134764, -0.0601188673523472, 
    -0.0457686770262082, -0.214787962347878, -0.0337068265079444, 
    0.0222578196965941, -0.182381900910112, -0.0200734302479084, 
    -0.0561639995226591, 0.0166750720703906, -0.217501058540153, 
    0.00298879765011355, -0.0785217245601355, -0.0112665114506351, 
    -0.169905684747602, -0.015596744462353, -0.0551812472604439, 
    0.0590029900136073, -0.227646110918767, 0.0350668051929911, 
    -0.00308491539965362, 0.00525052307360331, -0.00801571327495951, 
    0.00164801605007987, -0.0076366957352297, 0.00868685695467698, 
    0.0338283328870292, 0.032375887244845, -0.0452196563880689, 
    -0.125828255329775, 0.288696700392567, 0.219391991754963, 
    0.0344222560008892, 0.0444745062159789, 0.382556719840633, 
    0.193892188105178, -0.00545572156953279, -0.153131085709309, 
    -0.0890545750859498, -0.196225444427807, 0.948730259639177, 
    0.205967947781203, -0.0894712825962431, -0.51590228077489, 
    0.0226247005465195, 0.93223221600231, 0.565037546621602, 
    0.385562220460663, 0.811765486431841, 0.05724357862041, 
    -0.0807288239204031, -0.0501496320219944, -0.13204201024699, 
    -0.0503121939211996, 0.181476327255963, -0.0454210052585659, 
    -0.132747517639027, 0.0272812466575777, 0.0889015252124609, 
    -0.132362596144732, -0.0686702677418765, -0.121211400417386, 
    -0.091167948775678, -0.103837700120707, -0.0937121738782888, 
    -0.0441745824635427, -0.155050455516383, -0.00770120971781529, 
    -0.149226789282982, -0.0101676510578309, 0.00634556402748689, 
    0.0333831883707587, 0.00371717193446493, 0.0378780957652287, 
    0.0304943313142933, 0.0633959221488765, 0.0105797610192769, 
    0.0509711494565727, 0.031953999360443, 0.0651276516822329, 
    0.0388274056777896, 0.0520349332087577, 0.0381910621673659, 
    0.05158647183387, 0.0316611410665672, 0.0478165100319097, 
    0.0488066074915228, 0.0548468518758191, -0.00715796933483662, 
    0.0579858641699826, 0.0920901610714115, 0.123717072066832, 
    0.151780118651935, 0.0997828842614453, 0.0635456936343189, 
    0.13356509368499, 0.343151283095851, 0.243747281429898, 
    -0.121685471760406, 0.465651294418851, 0.383691360726666, 
    -0.086895333797985, 0.815187513605987, 0.430661587111026, 
    0.0578570191925391, 0.222256459364429, 0.0410455133076565, 
    0.542164940939457, 1.02140129580847, 0.307778311193723, 
    0.023141990440469, -0.00756949137575425, -0.00166746366558024, 
    0.0333303991900863, 0.00165429643177091, -0.0571860064832029, 
    0.0741265557949099, 0.0338327196491262, -0.0211105798202643, 
    -0.037439307955099, 0.00843740871844877, -0.113513175516112, 
    -0.0155247793055323, -0.0497619001395343, -0.0819701656898297, 
    0.0275960374572871, -0.0727323598548633, -0.0306087353431821, 
    -0.00860502126094445, 0.00411131877114477, -0.00407865710730813, 
    0.126595157553741, 0.21481864044902, 0.119798856242783, 
    0.0389784235691796, 0.0491081264638578, 0.118202785980069, 
    -0.125373581378421, 0.318976616905069, 0.453640537701169, 
    0.0350553822564504, 0.0227253246428973, -0.157159566088977, 
    0.673638903648063, 0.140091114015978, -0.0205766414501569, 
    1.32675071889673, 0.297456634751838, -0.0215551494152957, 
    -0.121738467230472, -0.234782322317175, 0.193358508611155, 
    -0.185977642119882, 0.176554420872462, -0.227140198887524, 
    0.118753744862213, -0.169524858401983, 0.11270387753914, 
    -0.0984997214373063, 0.233521257394181, 0.0323798842076159, 
    0.029655898491555, 0.15721145608833, 0.115338437084734, 
    0.0568688557965086, 0.0977119245079732, 0.119137150884538, 
    0.0996898193674285, 0.0397752837481339, 0.0306809258886771, 
    0.0460036817276364, 0.070109446938641, 0.0585265885099205, 
    0.0625747161215037, 0.044520155462357, 0.0539079064179076, 
    0.062883387400735, 0.0561155204951921, -0.00148626991110404, 
    0.0120714915117333, -0.104549566983842, -0.00896281566845983, 
    -0.0453819962562265, -0.048454726842727, 0.0432468342168531, 
    -0.119400759641479, 0.0618938541639758, 0.158815514179771, 
    -0.156513082411198, -0.00226060840793386, -0.189191477377252, 
    0.605461725507912, 0.29150743968485, 0.0651374902224111, 
    0.532045391076229, 0.363989513571487, -0.371734027545156, 
    0.49163026568852, 0.512565485700154, 0.150546062301799, 
    0.136232719163574, 0.0250076774919241, 0.619890445662758, 
    0.192415868357607, 0.185378504605292, -0.191005655874837, 
    0.361669602433588, 0.313720660753388, -0.056213349848702, 
    -0.201549488995029, -0.155813154161045, 0.0572989115471816, 
    -0.103747678339304, 0.0657825609094297, -0.238855093654496, 
    -0.00552317094161371, -0.119673043120143, 0.0538100342220431, 
    -0.132252613253362, 0.344929496351229, -0.0015708989175458, 
    0.340776576929665, 0.560706381192984, 0.171231333320256, 
    0.0451804315458086, -0.170304841293845, -0.00648885483491232, 
    0.480075002061315, 0.374734604478409, 0.19668781284948, 
    0.257235137865503, 0.335997340135681, 0.144182729374205, 
    -0.162113018113037, 0.562057376471328, 0.588267118254579, 
    0.177835737278177, -0.00698762641218885, 0.456685880985896, 
    0.420286307871971, 0.199847522572484, 0.112126658444476, 
    0.103848379266645, 0.109311816747709, 0.0760614470206425, 
    0.0820198810809018, 0.196190858726436, 0.102418472321736, 
    -0.128271934770122, 0.09051939957766, 0.39720492768264, 0.09412749301316, 
    -0.0991927345317827, -0.011886532737297, 0.418758714166548, 
    0.221256913524786, 0.122846459341738, 0.150391588302324, 
    -0.179237156128701, 0.470112071712697, 0.286873028579379, 
    0.114675226509894, 0.073957568989024, 0.0840331152363889, 
    -0.0558351211496006, 0.261864589250805, 0.308702591477552, 
    0.730772625832626, 0.497721364946056,
  0.285653508478233, 0.478306240889803, 0.0145669834921461, 
    0.0619869772657506, 0.0871647934012598, 0.773823461914334, 
    0.724260059703387, -0.0173886633149367, -0.152097033711608, 
    0.317534471263574, -0.0929215597605707, 0.538146372124093, 
    0.154427781121105, -0.220021473156197, 0.170857990779336, 
    0.576271014983046, -0.0398696542095788, 0.338371000612145, 
    0.7346555234998, -0.0732634199955393, -0.100563432896733, 
    -0.0672893870810891, -0.0602886027593858, -0.0805354333318466, 
    -0.0518658361848728, -0.0722744216183264, -0.0590284100551427, 
    0.0319060990124038, 0.215409001019802, -0.211380849813814, 
    0.178614694050549, 0.301571891318199, 0.163191558140306, 
    0.198636212739834, 0.195103954802628, -0.15443186116545, 
    0.55765553880778, 0.491198912511984, 0.0438206539776443, 
    -0.17060204849167, 0.142764269226418, 0.00828139489781014, 
    0.346297982912651, 0.72704649738101, 0.434839679116839, 
    0.146063088159592, -0.503158485467154, 0.037628361508247, 
    0.560053714651764, 0.201155143518913, -0.0702003223238365, 
    0.148893490149751, -0.165155621244072, 0.0853828733627312, 
    -0.390426187421108, -0.0740522294476052, -0.117344930389652, 
    -0.179748849698531, 0.18664830984599, -0.297812644292706, 
    0.0230547094190234, 0.102339327454186, 0.134469201771215, 
    0.136517680528287, 0.138654142305726, 0.110402418913657, 
    0.117279911385757, 0.157166353244335, 0.14431597943367, 
    0.0879702171222183, 0.133211610958373, 0.141547108794452, 
    0.149471782108112, 0.239268574625526, 0.242879297670872, 
    0.143922989111505, 0.180517216078325, 0.302944801041728, 
    -0.116154655551872, 0.121292580634084, 0.821066490656868, 
    0.354686656176288, 0.115792490533631, -0.172181313174067, 
    -0.118676912168882, 0.225739425955693, 0.440737045492288, 
    0.532808436194885, 0.439868766376607, 0.251301234713243, 
    0.0996439925472973, 0.0281498170360248, -0.117027746608029, 
    -0.111344010729408, -0.112413673541144, -0.245538082447754, 
    -0.106211533521733, -0.137922439513521, -0.176855073009335, 
    -0.0198639576950086, 0.00538507796975139, -0.166446561180489, 
    0.0705980596916318, -0.111539674737241, 0.0564629539111706, 
    -0.0741260975642182, 0.112735959331288, -0.191827455518711, 
    0.0417736744847131, -0.325534865792759, -0.125100416009314, 
    -0.0243294458284623, -0.00699930696252579, -0.0444995048356317, 
    -0.0918988711810577, 0.0503304186435503, -0.0109776158028738, 
    0.241431166315202, -0.0623377336172632, -0.244078915826837, 
    -0.225881111532561, 0.111477501242983, 0.313780980842097, 
    0.593914178321244, 0.500397232172241, 0.0982655984106376, 
    -0.576247524133557, 0.142202341712275, 0.6119297190296, 
    0.149350466186836, 0.117774570782832, -0.318074332763465, 
    0.429056084118122, 0.46409891609401, 0.210509666096757, 
    -0.198753088940986, 0.449813813649389, 0.42778513449248, 
    0.162208636568177, 0.101456725365435, 0.332938938978288, 
    0.229827268516445, 0.0684651103361235, 0.0601049884357105, 
    -0.0673779569103964, 0.314170920476602, 0.00849201294460054, 
    -0.0584167322933287, -0.0369318554727535, 0.23332333525002, 
    0.0904638591617411, 0.148667723972926, 0.297444476575514, 
    0.105325042503601, 0.0504049675417421, 0.153667569717066, 
    0.488785053483665, 0.181883687614383, -0.00749840673399807, 
    0.0932652105536841, -0.139831688567332, 0.101442072562331, 
    -0.121902821400816, 0.090494384631587, -0.0693115371710534, 
    0.0981349313558006, -0.115077960876827, 0.056088631215184, 
    -0.19214820318727, -0.050733512432559, -0.00796620345249501, 
    0.056693053675231, 0.027099505119414, 0.023484333372177, 
    -0.0256219317482441, -0.00765789838410533, 0.0290934326430654, 
    0.046079786527911, 0.107839897216856, 0.0167298122270562, 
    0.0705581944279465, 0.0972154892893108, 0.100982064190383, 
    0.128181916979879, 0.141192819723984, 0.109130591718926, 
    0.109964648889941, 0.181029913841873, 0.126400569352144, 
    0.00464311336195673, 0.134151706027247, 0.273085284373061, 
    0.142478357874756, 0.185991440255237, 0.397029337948483, 
    0.164804594504738, 0.160279570068668, 0.62633747451887, 
    0.244758779231256, 0.0255576924912502, 0.035834201445395, 
    -0.352831236736933, 0.332059575120791, 0.578780547322341, 
    -0.0200623775842706, -0.0331377980084136, -0.329477679324744, 
    0.180324438414144, 0.538349354826926, 0.169050699268151, 
    -0.107269199522018, 0.109458160853578, 0.132399996897257, 
    0.0235925650200957, -0.0128773445507127, 0.00747322824908336, 
    0.320636561630086, 0.0228296239706117, 0.0176784982970477, 
    -0.0120234304582463, -0.0515593706973366, -0.169194253937289, 
    0.0938936565639947, -0.15280648464064, 0.00331005245068382, 
    -0.0931535957990581, 0.0305591613694353, -0.113048117294813, 
    0.034940400242828, -0.237424790282967, -0.0358481860129831, 
    0.0439098198656331, 0.124955444853715, 0.155810348269054, 
    0.120441654753252, 0.0901020523261693, 0.16579906126435, 
    0.215508661340581, 0.150728553586279, 0.106060005323623, 
    0.160927122943448, 0.142041361740929, 0.286107559661199, 
    0.35787046984143, 0.179460206699937, 0.112952626557127, 
    0.460107656176414, 0.411133910911388, 0.223388625254214, 
    -0.0363803118932474, 0.782412107203341, 0.046881547432575, 
    -0.265001206918858, 0.101334623567703, 0.764316883166494, 
    -0.236105136491803, -0.364647092358732, -0.0978937547766949, 
    0.805451356588116, -0.0386877752350859, -0.0661028865879314, 
    -0.151540852826474, -0.0724308835844568, 0.288503241229028, 
    0.372814334561061, 0.11817411771137, 0.035576292265053, 
    0.951757532207101, 0.12021320078084, -0.0210513999677487, 
    -0.0482452096935342, -0.180098115352837, 0.111694666867336, 
    -0.414308393213154, -0.0131290932131044, -0.214116779743438, 
    -0.0528490552459187, -0.155306911031391, 0.235846367112424, 
    -0.144652823127341, 0.289073796303522, 0.10458254929701, 
    0.405398818917232, 0.466014124851063, -0.0134672214907939, 
    0.379875992297935, 0.714173750711414, 0.174030204650555, 
    0.138504162999219, -0.262546072643449, 0.159142190936788, 
    0.449303097618597, 0.195171639475036, 0.143234128319392, 
    0.555670306147216, 0.169977050784617, -0.0389016770130954, 
    0.170914735372068, 0.434379962125778, -0.00821566391258895, 
    -0.104969668060488, -0.108034396910537, -0.000932505589388899, 
    -0.0837505246293842, 0.00791133535651999, -0.137823198488019, 
    -0.00377051065432324, -0.0757433974000652, 0.00633123954313594, 
    -0.135835772676433, -0.0619578041931647, 0.200267698919143, 
    0.115638092129363, 0.0249139221078081, 0.116849294187547, 
    0.128459298543849, 0.342115516727576, 0.27000198172162, 
    -0.00183083860705588, 0.0433991157551673, 0.432601798347443, 
    -0.225211211186151, 0.25950529678672, 0.402558314554346, 
    0.378552722684825, 0.675204578942668, 0.405099226465666, 
    0.0279697683074362, 0.94937625434204, 0.331072471174111, 
    -0.0541207313394191, -0.00798043360149432, -0.0847946295170833, 
    -0.00771921592568489, -0.0800110175223536, 0.0744728256559266, 
    0.0422610005241849, -0.0957051490010108, -0.149869564954287, 
    -0.155990769758036, -0.132441157488701, -0.105220893121425, 
    -0.0367775224544845, -0.147944624769922, 0.0533309634036748, 
    -0.139103375764531, 0.0508312164032426, -0.117861809873768, 
    0.0416213434869361, -0.141910318439965, -0.0043717658857531, 
    0.0282518882692915, 0.102939558051003, 0.114397786173404, 
    0.09301899904265, 0.0918536099612056, -0.088358798151685, 
    0.493701753906908, 0.187919278265004, -0.366631179453528,
  0.297794969662477, 0.357574219248014, 0.318811588710128, 0.4637053481174, 
    0.298751074254106, 0.0416610648557398, 0.251811129027464, 
    0.42041070460184, 0.224888038851876, 0.105479256416885, 
    -0.0836145861849371, -0.169588653874681, 0.302602756863006, 
    0.456885490804821, 0.19155138323113, -0.165800747123769, 
    0.272169239750218, 0.31757248633617, 0.148023560790119, 
    0.339755987247224, 0.2211450992763, -0.111326590195631, 
    -0.105770595188054, -0.0152601136043422, 0.219722081946032, 
    -0.0795705672800552, -0.246936306149147, 0.025328383085416, 
    0.220429650523493, -0.0409903083534193, -0.0806800163893155, 
    -0.164060597503497, 0.17478194810242, -0.221992721858974, 
    0.0854247831248534, -0.33349794535893, -0.0255723074022509, 
    -0.15076735514338, 0.0383447301886799, -0.344434120011536, 
    -0.0294455124326678, 0.0693206443570795, 0.082017664368681, 
    0.181439563500685, 0.212806483168787, 0.142501525927556, 
    0.115948301980018, 0.189650810423337, 0.196424940828975, 
    0.14270081196789, 0.178173963254489, 0.206449044393959, 
    0.286207108565951, 0.268897692254871, 0.135787351640563, 
    0.213428258789318, 0.510648379274555, 0.238669237616614, 
    0.00947627222111672, -0.123623293338265, 0.392327398488784, 
    0.556185805450937, 0.0913462055843154, -0.241024637695228, 
    -0.0525788042576227, 0.552504306591766, 0.0874714028464426, 
    0.00559035072498673, -0.0180418966555635, 0.54431117902938, 
    0.116833046225763, 0.0863714181757193, -0.0651795530477119, 
    0.273255301240615, 0.0678433696794516, 0.0723222562833244, 
    0.200970547270306, -0.213272024630173, -0.0883790265957885, 
    -0.0810938997238419, 0.0532496804337264, -0.251333459573048, 
    0.1275565727927, -0.128286088592614, 0.043650413357633, 
    -0.222214121482233, 0.017565796055795, -0.157254211671826, 
    0.0376328820016758, -0.337849272669415, -0.0548651694900625, 
    0.0320490006126933, -0.00780445692809977, 0.0508478336004322, 
    0.0924595153585153, 0.056811218364412, 0.152365498163255, 
    0.136686020613175, -0.181576937616112, 0.117963351344384, 
    0.45285655782044, 0.231881855696907, 0.143470396785309, 
    0.619975069266047, 0.266745585916581, -0.195981735886619, 
    0.145309374298381, 0.0229069212860881, -0.0823820915110868, 
    1.16551385866598, 0.57821009140071, 0.0873068841916278, 
    -0.0125636211695498, 0.087610456873997, 0.186155745528282, 
    0.0912217410827235, 0.079446929518208, 0.575873445349024, 
    0.23191023834353, -0.0120488229344849, -0.0490436298870019, 
    0.132377642945663, -0.260983242097265, 0.0474418367662256, 
    -0.3300222807487, -0.224021273168369, 0.0490486330905273, 
    -0.0816559161453094, 0.252031405107434, -0.144322378550921, 
    0.247158783005614, 0.206606857171241, 0.0499202561183747, 
    -0.125343842679488, -0.0596720385308668, 0.512736360048061, 
    0.122204245671315, -0.116308202005341, 0.138459752320367, 
    0.402475422152607, 0.130532957496822, -0.351634479552479, 
    0.266479522794012, 0.671442950833644, 0.155088295217107, 
    0.0118369380561132, -0.207758375052003, 0.0123789179390602, 
    0.516393954003567, 0.429609638656311, 0.203818851468767, 
    0.197883701285714, 0.198200285168383, 0.245277269925566, 
    0.307869625153075, 0.2209503088987, 0.126064761558818, 0.189639630685953, 
    0.219832418172188, 0.0561634111900387, 0.0743089226475205, 
    0.518527213116536, 0.173556196372193, -0.0950393981446335, 
    0.174073183069504, 0.462345976973692, 0.0264146902620432, 
    0.096866748668039, -0.116370699055649, 0.102007388279643, 
    0.366795688890976, 0.274425545276203, 0.00546642701282819, 
    -0.139117223922501, 0.110671504019246, -0.328168832214994, 
    0.437978585299294, 0.454358125014263, 0.222001616451702, 
    0.132344765530828, -0.149458383626683, 0.118453704530101, 
    -0.234748007546029, 0.044229486621596, -0.342254026724964, 
    -0.121653422402694, -0.0793542857935602, -0.209757835206403, 
    0.12176486589856, -0.199191199962924, 0.0966980648791489, 
    0.0328191015239511, 0.0696218660551973, 0.0497517637896487, 
    0.0809676425450362, 0.0208185738279447, 0.0622687696887089, 
    0.0694348661277481, 0.0741937715021956, -0.0192935051364427, 
    0.0559718472249976, 0.0753797492976264, 0.090383544819092, 
    0.182578545658996, 0.166375761645652, 0.0632271504274021, 
    0.0404904884147944, 0.333017917904709, 0.182667166328769, 
    -0.151485941129958, 0.358488940682087, 0.346565722736065, 
    0.0473457277558068, 0.10023852899333, -0.350751498852324, 
    0.130298438615526, 0.559125741208085, 0.172442388332893, 
    -0.120865026173323, 0.0700568944620709, 0.286785969265351, 
    0.386925487585955, 0.178243108144932, -0.0561226847925788, 
    0.0449729052101535, 0.0755858862887616, 0.610622998730797, 
    0.179107830505392, -0.24485840820415, -0.0836705391595462, 
    -0.24515946167904, -0.0440996773042153, -0.303636228782997, 
    -0.0772157598103252, -0.258666002121864, -0.114270216751988, 
    -0.23839876608712, -0.106974150336455, -0.192365977045472, 
    -0.151446486770932, 0.000326782731000855, 0.0201542250174052, 
    0.0222588222498217, -0.00760671745587133, 0.111016926853768, 
    0.0165296036128889, 0.0523930530165647, 0.0379058176878072, 
    0.0345673764980509, -0.00705405042114508, -0.00199558290152961, 
    0.142684977744989, 0.132823030267839, 0.0376852826797663, 
    0.0523083844217018, 0.263591454450811, 0.146145179880657, 
    0.0853077162551272, 0.19649766072592, -0.166214227854985, 
    0.53296563776731, 0.343107167794327, -0.00810593762408005, 
    -0.117891578789879, -0.0219808058164783, 0.632087985406369, 
    0.36872709430681, 0.204673053885342, 0.800944324175393, 
    0.442949001703079, 0.0581607655277924, 0.0585661480984545, 
    -0.082524004743582, 0.0807832988582803, -0.0137794696239643, 
    -0.039526966583641, -0.0154219415732842, 0.0108075763476899, 
    -0.121306146582194, -0.19659086976591, -0.180636810041866, 
    -0.0169537204076687, -0.150136406841717, -3.45576430858391e-05, 
    -0.0638095162985524, 0.0381466748948385, -0.3851494135244, 
    -0.0442709680505299, -0.0572526324725077, -0.222360145778818, 
    0.057718440074758, 0.0227852572824901, 0.0250730441262552, 
    0.209805452459115, 0.164984854873608, 0.0378929430240416, 
    -0.115991858921351, -0.0134667500722858, 0.408853292543277, 
    0.184698263638933, -0.132718434520478, 0.0928225287399083, 
    0.394576398952474, 0.771402143251748, 0.409946897076542, 
    -0.227176262321865, 0.475326428753957, 0.397312201462556, 
    -0.00649851695660467, -0.0269940302711541, 0.578434722489208, 
    0.510039525284357, 0.108871403426815, -0.220458206694083, 
    0.0917365504510658, 0.519651354570699, -0.0174867022391472, 
    0.00203313237331708, 0.915460351858873, 0.0356100291731713, 
    -0.173691327536731, -0.178736662001536, -0.122540627265138, 
    0.153234547708817, -0.103705797476739, -0.213843970605111, 
    -0.0124148248555535, 0.0978714395060828, -0.105532699835569, 
    -0.0511510692319507, -0.0555309113328776, -0.123636718030162, 
    0.0333129124084128, -0.0468233834087897, 0.0229867558611632, 
    -0.062163175736261, 0.0454086244932227, -0.0563187136358764, 
    0.104869221226709, -0.055914942931413, 0.229612282034976, 
    -0.102236764750717, 0.526900742813811, 0.458344195995921, 
    0.0619620920756233, 0.0187706399193175, -0.258218852763382, 
    0.207575448018825, 0.46283099576836, 0.265259757615224, 
    0.157037229913921, -0.159976601826031, 0.379123856546132, 
    0.449593949378574, 0.137183415827768, -0.301477251755133, 
    0.210431536312698, 0.614399487903014, 0.26290358341154, 0.0914365188928355,
  -0.0230571504554317, 0.0750029165615763, 0.11698536459414, 
    0.129340809419697, 0.16768755503714, 0.270192138164176, 
    0.245012817339708, 0.161740867474887, 0.173911524205518, 
    0.209893830537667, 0.237085361434623, 0.245766134925472, 
    0.250352140301052, 0.215421485414181, 0.126472969461312, 
    0.19608362744536, 0.36721171273003, 0.161807995761509, 
    0.0104714192804241, 0.0318216166041466, -0.0766585274306181, 
    -0.365168540009685, 1.06916506325234, 0.328047394347339, 
    0.0535054605301483, -0.0453616060821563, -0.108266002690829, 
    0.74586915105602, 0.173008401140945, -0.0520557044378503, 
    0.505935231659252, 0.263977950973087, 0.0384820155429637, 
    0.00503723412029219, 0.0111527710828317, 0.0139999649307915, 
    0.0237967704766805, 0.0273999725689355, 0.0168557829825564, 
    0.029314924709143, 0.0476282541062764, 0.0364544817151975, 
    0.0209081652481266, 0.0211581970883316, -0.0116130798887118, 
    0.015675318977939, 0.0125311998964223, 0.0328752855261642, 
    0.0451298077198788, -0.0145448960988209, 0.0685664600491274, 
    0.0971097862521123, 0.121408111548538, 0.156934206838954, 
    0.171036654874399, 0.157678654976012, 0.167649853636349, 
    0.198072524643435, 0.178419978858423, 0.175385515906823, 
    0.244494439405347, 0.174933304483496, 0.0755056649521913, 
    0.302573557545833, 0.416304936894174, 0.184451159544532, 
    -0.013708545208827, 0.325421278481339, 0.44896564851212, 
    0.148059500112654, -0.0121150724973458, 0.107267524956797, 
    0.333443589590717, 0.187480003776163, 0.204838584699114, 
    0.607140413967907, 0.617760779928672, 0.291208984729171, 
    -0.163970958170522, 0.811842777249507, 0.333888065364297, 
    -0.0048322824963881, 0.00930517141545348, -0.0124001355536061, 
    0.0269471254041556, -0.104008393401167, 0.957742722239256, 
    0.0968226508515338, -0.703363238395025, -0.305535684834218, 
    -0.264636069006019, -0.22375687942752, -0.140797050579584, 
    -0.358388741651026, -0.031236216401679, -0.466393769781335, 
    -0.166106661305183, -0.248423351596278, -0.294305454492566, 
    -0.125399156550655, -0.046345990030674, 0.0387772902489629, 
    -0.0199413585680262, 0.0613082675105949, 0.00815082559200794, 
    0.08914999342461, 0.0228035826065294, 0.0731466490122405, 
    -0.0179677696095516, 0.0440168439968649, 0.25229380956635, 
    -0.0243410654630713, 0.0861907895676867, 0.4375233516643, 
    0.335553017602599, 0.0963675742297804, -0.00531985149928532, 
    -0.110435052949125, 0.483282426720563, 0.0481654223515418, 
    -0.108281463987611, -0.297266743066995, 0.630596128906543, 
    0.599464191037169, 0.274092674837765, -0.406994798999096, 
    0.338489551666174, 0.580158255978795, 0.0976866875311827, 
    -0.188629346960925, 0.0878508993510672, 0.72353567569996, 
    0.034741862654836, -0.110194058880205, -0.0741606625456748, 
    0.574398618675785, 0.267363475102822, 0.229085774563107, 
    -0.0445150610604662, 0.504260523719233, 0.212685376761732, 
    0.029915128892065, -0.0230099303646938, -0.159367130007177, 
    0.0536767461506926, 0.19450074790922, 0.0545176394102169, 
    -0.072757058601407, 0.166099061589598, 0.416325988840877, 
    0.114810686410994, -0.0746097309080923, -0.153584332030003, 
    -0.0337982499479804, -0.0922077512108891, -0.0658589147882277, 
    -0.0470334215269092, -0.0970018864204813, -0.00665162258061203, 
    -0.114243174956002, 0.0151328331806554, 0.0680413860217054, 
    0.064310456427689, 0.189971385105761, 0.199899050217502, 
    0.0737888821425249, 0.071603625813992, 0.222017972016098, 
    0.23600890525614, 0.103169830407897, 0.255365069800124, 
    0.817318903073164, 0.268108183709702, 0.0416275818862098, 
    -0.025888601199292, -0.437785508343984, 0.841261029759331, 
    0.364820288316909, -0.119750122891133, 0.413907934536444, 
    0.489274332782245, 0.191593795145316, 0.128843781381725, 
    0.0847618543178019, 0.400874837184672, 0.147500811223583, 
    0.199716795157607, -0.542230335168372, 0.456189554046903, 
    -0.0650775109617963, -0.317485728039039, 0.166321677127087, 
    -0.291794921790636, -0.0267309615412707, -0.27560940481468, 
    -0.115649093967302, -0.156230236486459, -0.191003906671862, 
    0.0599506222486436, -0.227470155556535, 0.229034647913571, 
    -0.0679831637695504, 0.0668886721609028, 0.494559713522731, 
    0.14629689665262, -0.00186300857877007, 0.165242891191249, 
    0.279473735366078, -0.211961260977141, 0.517423035554124, 
    0.596338398587222, 0.151253350404769, -0.143238717980553, 
    0.60799515562145, 0.469418993072555, 0.172876403942352, 
    0.069892343232712, -0.215861362162612, 0.270903015418934, 
    0.560116106541306, 0.234990690981625, 0.132565907801459, 
    0.266538803296978, 0.29075931805754, 0.155897874419551, 
    0.196169699026047, 0.371951488031628, 0.225094382455467, 
    0.0878025810965088, -0.153914218557749, 0.275505185292706, 
    0.400234978365616, 0.181449803123497, -0.196533873477998, 
    0.277850572610779, 0.374110542045692, 0.0769528785765504, 
    0.0642060631322577, -0.25531738931646, 0.334585129979615, 
    0.335739121925331, 0.0347180167962671, -0.0515019644497735, 
    -0.0696281361518103, 0.45296659233638, -0.0209892424847138, 
    -0.0578339640858321, -0.124556856844809, 0.39653649094872, 
    0.0740361157049456, -0.0926354475071788, 0.0370502130998385, 
    -0.047341955707329, 0.0617772238699973, -0.109495935561603, 
    0.069188269707555, -0.336441402369254, -0.0494684037329565, 
    -0.143642352968584, -0.153101818450702, -0.0281018455090273, 
    0.0851840372640798, 0.121113986338607, 0.119604981240626, 
    0.151487666524286, 0.156898282232417, 0.16043894777188, 
    0.199323735260451, 0.168783605861348, 0.0862118855269142, 
    0.0573545343228078, 0.284881075139543, 0.350958940976752, 
    0.150303983750818, 0.021143392563045, 0.39577017244684, 
    0.351798190945371, 0.136752713484431, 0.409047244091368, 
    0.40889015160449, -0.0140250217011921, -0.0461955228022166, 
    -0.208378549851372, -0.265031997562325, 0.734932777656874, 
    0.131253578181045, -0.00563654952201231, 0.41744599478677, 
    -0.250639588302707, -0.295281346215941, -0.104663759425865, 
    -0.250339421185573, -0.0758969756659001, -0.275737917794443, 
    -0.0048352976085717, -0.219402537242078, 0.0543147173589603, 
    -0.219182957413197, 0.0849512574373674, -0.284804199430082, 
    0.0132915259506556, 0.00678682696745406, 0.100190619000832, 
    0.0101263426271287, 0.113864278003138, -0.0790887573899113, 
    0.022801378584658, -0.016723461880969, 0.0172045943534588, 
    -0.104865928853486, -0.0237632347313932, 0.0279287923920418, 
    0.0887055340476666, 0.0889508995742563, 0.0576576451686331, 
    0.0295549384224493, 0.0817136057352715, 0.136375533730908, 
    0.0779480259299211, 0.072648506416154, 0.20394520449714, 
    0.0335294422973975, 0.0314213658350048, 0.503795858632171, 
    0.265015364744525, 0.0836647695285136, 0.0309127800366051, 
    0.636718081807201, -0.0178532289686162, -0.0828762126275442, 
    -0.222905120567391, 0.269930657746108, 0.620966636832149, 
    0.269782363199379, -0.204064305789866, 0.272681473858625, 
    0.540877631644035, 0.178441417532323, -0.173489451316415, 
    0.339669980373615, 0.356859808640361, 0.120232892517241, 
    0.0685975038935135, -0.00401630401990354, 0.222021474578534, 
    -0.200786054951688, -0.169995793640937, -0.143013663085867, 
    0.0259379044831789, -0.0225935248999604, -0.1088433751643, 
    -0.309719246522536, -0.020322256464591, -0.141077962079475, 
    -0.041567739832009, -0.301675049026177, -0.0419374110543073, 
    -0.156862150438187, 0.00792587803644185, -0.350383590313033,
  -0.101910891857913, -0.0665644006017068, -0.0144743249224023, 
    -0.112775730602795, 0.14076384905119, -0.0561351627493589, 
    0.0549181835247067, -0.0772499678839888, 0.0163000537926085, 
    -0.161179048710006, 0.00443282036057335, 0.00127651469961392, 
    0.168734093890863, 0.193152274698375, 0.0758859685320351, 
    -0.0359150304033349, -0.00396843108935567, 0.290825914097152, 
    0.194935924675251, 0.0992363968206407, 0.387848331312399, 
    0.240752340368388, -0.123323591906165, 0.0374449292824805, 
    0.739425353543175, 0.191263697467289, -0.339523820445354, 
    0.407197264489633, 0.632082133364469, -0.0327223864802771, 
    -0.171665590004822, -0.159911596262709, 0.537378025346256, 
    0.325763525864572, 0.103210956036867, 0.054786408743063, 
    -0.226145564965001, 0.542774121724475, 0.346430268571562, 
    0.121053601538295, -0.187512973724522, 0.197118249187371, 
    0.298943942220829, 0.0110525939721798, 0.169714512532271, 
    0.509965480815387, 0.145958955181094, 0.18491173098461, 
    0.208608233140365, -0.194916787754546, -0.268256788777904, 
    -0.0150715259794556, -0.131030855464278, -0.0319903746674683, 
    -0.117658102004219, -0.111526701443274, -0.133558884579644, 
    -0.252718684431311, -0.0257932798192346, -0.214151458173336, 
    -0.101791772306069, -0.0295109783578926, -0.137934869226607, 
    0.0859735760011329, -0.0488228837956042, 0.0727320140393542, 
    -0.11588398430259, 0.00443213953555224, -0.222476198135296, 
    -0.0799829368542404, -0.00840826091473412, 0.0274296397734355, 
    0.0446433346588539, 0.0542931393194826, 0.0526033621627559, 
    0.0440048035938665, 0.0125610996500783, 0.0465731150873107, 
    0.0767871393851926, -0.0438204847699957, 0.192783613307101, 
    0.229889921931443, -0.0418120078590129, 0.365332578567643, 
    0.335048629309236, 0.0652919344474969, 0.398269532433134, 
    0.444462377433435, 0.102837640690998, -0.059871041847795, 
    0.0589607290249453, 0.11156354981452, 1.14207399004433, 
    0.370152585259892, 0.088072825977695, 0.235252234391104, 
    -0.0788547251062254, -0.0623831961194876, 0.310528796650815, 
    0.764797479749901, 0.0942244361626071, -0.141658508181222, 
    -0.109334780097758, -0.0823857124584134, -0.117592375419852, 
    -0.0285575123099364, -0.128351281328709, -0.061530361808662, 
    -0.0972596345836448, -0.283388372553949, 0.130265942332192, 
    -0.121077863180085, 0.0877367303432013, -0.0367656177116545, 
    0.130517148177674, -0.184935035022937, 0.0822534383684935, 
    -0.212472084063166, -0.0412290023421184, -0.0962350233607249, 
    -0.0129751981480032, 0.0477192214729962, 0.018408874734417, 
    0.0439624606954837, 0.0235192665634829, 0.0504989063970377, 
    0.0279431688739165, 0.0496572922731844, 0.0183668003592993, 
    0.00291660344040556, 0.0659829676957217, 0.107405043952144, 
    0.125849900008581, 0.136308604737084, 0.147084264398713, 
    0.125929793159291, 0.12486120064239, 0.180292323576637, 
    0.152073536317671, 0.0718441379649246, 0.128231577578316, 
    0.247666754044625, 0.205842534074915, 0.11265636894329, 
    0.281983614461783, 0.3936824023936, 0.182366522751495, 
    -0.0564558099879355, 0.323345171991901, 0.490069884594166, 
    0.188149056089073, 0.104849576877322, -0.262537433522544, 
    0.169877405036496, 0.388355372496509, 0.557091191010797, 
    0.231901510875402, -0.146624516409721, 0.0333671390332351, 
    0.635305267968237, 0.0156767103001385, 0.0403846793938833, 
    -0.0964184094593444, 0.200365004455222, 0.182147700393183, 
    -0.0835204568918907, 0.0791201793930788, -0.129611863981092, 
    0.245224240133876, 0.11613627238747, -0.0766441361879203, 
    0.0169744446927457, -0.0937461169561413, 0.0357324946110075, 
    -0.192978711009642, -0.0026612805159328, -0.341654608680659, 
    -0.145577980786677, -0.0412262016554156, -0.234587923902711, 
    -0.0231667473373469, 0.0753636384154957, 0.104961342388361, 
    0.119155952893288, 0.165597053042796, 0.206254613837744, 
    0.202512681538256, 0.127312742176879, 0.020446490499279, 
    0.323915727238731, 0.394020669435263, 0.118340731999585, 
    -0.187592223818849, 0.399226188714347, 0.513868410842161, 
    0.177172452598337, 0.0358464935782021, -0.13819705023299, 
    0.145474946105503, 0.501543283749016, 0.509019160655176, 
    0.270210375237186, -0.118556550109395, 0.719783081283409, 
    0.290565657742748, -0.134852270266473, -0.26897798891233, 
    -0.177282355975663, 0.589939618385439, 0.101946199227789, 
    -0.0625107467226838, 0.06864695793217, -0.262551404762215, 
    0.00689504401106134, -0.295215669898069, -0.197957268916085, 
    0.0362706571569623, -0.124376436168526, 0.133683300331716, 
    -0.219916069773922, 0.0278713442763065, 0.109619720363783, 
    0.128445634176592, 0.147477188450961, 0.154151214545741, 
    0.131092444951802, 0.140203112910954, 0.189054638922756, 
    0.157793674629661, 0.0901135366573839, 0.186266851775321, 
    0.219555700665679, 0.160796450704396, 0.168660181304598, 
    0.273251891423667, 0.361411597585375, 0.247408974500227, 
    0.0676498326345923, 0.0073338288153495, 0.387640314514473, 
    0.583522948140779, 0.184857847119743, -0.183873620105409, 
    0.145681804842782, 0.313185023375985, 0.192168310638779, 
    0.673723586750559, 0.452041909634122, 0.0920511963341695, 
    0.51854577407765, 0.256092811670015, -0.12686547892119, 
    -0.0855748387011219, -0.12466380748579, -0.0552113004385919, 
    -0.0734964042752087, -0.139493964904857, -0.100386017524941, 
    -0.0770926208236564, -0.0956190173038396, 0.017573007009746, 
    -0.0963518176641797, 0.0449534672427562, -0.0673945069317027, 
    0.0207084430120172, -0.0794789102075811, 0.0264605495884803, 
    -0.0507506594805417, 0.0337155115891579, -0.151723438649973, 
    -0.0173190833094474, 0.0560377725293809, 0.01702364560113, 
    0.110608971691911, 0.127954463916372, 0.0545749188964413, 
    -0.00338556679513913, 0.304128047333508, -0.0673368839575486, 
    -0.0841068835346809, -0.268088592361861, 0.545379990125785, 
    0.275429794244544, 0.13701952846134, 0.242702288167421, 
    0.00933686187898379, 0.959842067823808, 0.19107564659078, 
    -0.040381215271299, -0.0518353304716729, 0.255835844429125, 
    0.556319457802146, 0.302815094048434, -0.0736953701011588, 
    0.289437899509178, 0.225832547131032, 0.283362301458197, 
    0.479419984235205, 0.138610158151784, -4.86134017523981e-05, 
    -0.212852253044227, 0.0487071219581905, -0.173955880914851, 
    -0.00898476305402975, -0.278497559095863, -0.081862782126482, 
    -0.0485862993936493, -0.119020173125508, 0.222434508398059, 
    -0.221182842211849, 0.137954667323455, 0.193937186337038, 
    -0.117569294245476, 0.0993870598608771, 0.508036086039793, 
    0.147100300802689, 0.0934434640958093, -0.123961934614201, 
    0.569859199511539, 0.160982841075583, 0.0171778592561431, 
    0.228316080999714, 0.835178732959324, -0.0686552451532604, 
    0.172364225177373, -0.352217029025138, 0.831399054879596, 
    0.200320806945668, -0.229813554389042, 0.350970104512548, 
    0.514929945553308, 0.196363436224528, 0.149567906285262, 
    -0.236640640211309, 0.265389780999526, 0.356964088769421, 
    0.208979311043177, 0.133050076964427, 0.0718954863430528, 
    0.636126107727137, 0.055251492851129, -0.0906117739595043, 
    0.111439617534394, 0.322818877075932, -0.0399665646825507, 
    -0.0491737239355273, 0.44945799014096, 0.29989342850738, 
    0.197371614885839, 0.0860972669956257, -0.147446330735978, 
    -0.133670118258926, -0.264419041342904, -0.185146949385664, 
    -0.221170333794562, -0.188999943740285, -0.1655005139357, 
    -0.237180282494475, -0.0953822227181034, -0.216635715803483,
  0.0310012986670766, 0.0890634003433083, 0.114067230747023, 
    0.12767491971047, 0.192568678847066, 0.236596225163285, 
    0.163343603083478, 0.0473239295893946, -0.0249022969557223, 
    0.473903878143168, 0.305578008411671, 0.0245696472342068, 
    -0.160379601350703, -0.175197292346261, 0.596415896738811, 
    0.392132310920365, 0.155842962704443, 0.674130619863577, 
    0.278195587218669, -0.0364837367924678, 0.138030157931236, 
    0.534639690933789, 0.112509855210288, -0.0427726225419062, 
    -0.107442433989362, 0.153198008285355, 0.74537752652894, 
    0.236826195062857, -0.0955738358875088, 0.197340819922105, 
    0.375016506797676, -0.0463427421854773, -0.038376528642382, 
    -0.00814061749864557, 0.113049015682406, -0.163609692755822, 
    -0.0366815299749841, 0.0801024566385923, 0.101035740116053, 
    0.0915613005207871, 0.057381193453542, 0.0647664026640131, 
    -0.0680894905199458, 0.0347359162123602, -0.0917042395026489, 
    0.0433328754450632, -0.180691979481101, -0.0244939058256347, 
    -0.331456695545941, -0.136364446291718, -0.0257007300551302, 
    0.0719777457623573, 0.0647198427027794, 0.0676951742729176, 
    0.0840533843734591, 0.0812123066189639, 0.0454217323155419, 
    0.0803002299210137, 0.0610683465214057, -0.0141473449697309, 
    0.0871693741320734, 0.200328672919469, 0.135255840449808, 
    0.089777575827235, 0.326076700347829, 0.280158153922906, 
    0.0878399584139529, 0.0346138229591608, 0.477897169870351, 
    0.22425847501032, -0.168018286713478, 0.297506085223885, 
    0.595826201443235, 0.125091089682038, 0.0649535165395485, 
    -0.189012274494316, 0.615480124648523, 0.27225915776685, 
    0.0874039126990971, -0.160953629671249, 0.274168105606495, 
    0.392163422632804, 0.121315187992693, 0.0635277720511777, 
    -0.202656850461388, 0.181104162665612, 0.143981752678789, 
    0.453418642458032, 0.467862050381049, -0.0942047862634972, 
    -0.16976917077566, -0.185432171900762, -0.0378027352012538, 
    -0.0740222111368538, -0.137179299096344, -0.117320820531618, 
    -0.120106885936874, -0.0352377150325884, 0.00452383758374603, 
    -0.0122105893076665, -0.0355365288747983, 0.0415155887218021, 
    -0.045153323177977, 0.027573416675321, -0.104673191023428, 
    0.0212721972581255, -0.117401882259571, -0.0264976271450756, 
    -0.201959909958709, -0.0959791340246505, 0.00470440371422239, 
    0.0565615248957049, 0.0315521044947318, 0.0377405863515805, 
    0.0829130646375479, 0.0361490023853931, 0.0440396115254726, 
    0.069134631781046, 0.0653062780269786, -0.00845041070390543, 
    0.107018781417994, 0.159002152668873, 0.0868659050628703, 
    0.165435362321562, 0.315380848106843, 0.176028782239711, 
    0.0423200731244965, 0.181224329371097, 0.216031319950876, 
    0.0452569631884762, 0.649367279977486, 0.354152047242017, 
    -0.129412744942243, 0.248579821597824, 0.541268663130159, 
    0.142338418102362, 0.197838655693763, -0.133899698004009, 
    0.681494908373386, 0.190066641916548, -0.0226301025392004, 
    -0.0883245421678766, -0.112804256031042, 0.237452164283844, 
    0.23171281223776, 0.101226790462083, 0.294374943281795, 0.12116565855955, 
    -0.375852537099265, -0.223232718462819, -0.264782118859779, 
    -0.164958016270202, -0.240621695619328, -0.233745327528408, 
    -0.131127004895635, -0.241248890777532, -0.0273500482377892, 
    -0.19536884588134, 0.111069554961424, -0.242687817474323, 
    0.0878975617676021, 0.0304604498645884, 0.0582921321190653, 
    0.0223377592433259, 0.0384237509855244, 0.0372789041978046, 
    0.063524052450302, 0.0504680420890518, 0.0883918510447055, 
    0.0036665013347766, 0.109021672619926, 0.0849503483940696, 
    0.139351181246696, 0.235782756565142, 0.203260214279717, 
    0.0467019058093851, 0.113298023843098, 0.415362602281219, 
    0.300583210843682, 0.187110710152171, 0.161072352061276, 
    -0.196958911061206, 0.187596163679007, 0.328851166084313, 
    0.304842608601405, 0.303134753193698, 0.784632692794068, 
    0.511260334582964, -0.0946489142319704, -0.0844600810220644, 
    -0.0346789472984208, -0.262054834266426, 0.0717347774924493, 
    -0.234883739572313, -0.00150001643258996, -0.13817010585466, 
    0.0665104795831622, -0.246952539101391, 0.0692825306466089, 
    -0.169230332324198, 0.0815887274929795, -0.00353339640777824, 
    0.0843317686223135, -0.00250830231655579, 0.0744964073132246, 
    -0.0443465888214065, 0.0319489401938406, 0.0536752214424305, 
    0.0684910041332201, -0.107133741450953, 0.0203710235482258, 
    0.0719921283013679, 0.0630920001347424, 0.0817959158110664, 
    0.145089363283086, 0.122954503224906, 0.0499683540278329, 
    0.00609361048938349, 0.390716483126493, 0.143389495385103, 
    -0.136845104290458, 0.0930026367583115, 0.583435214359945, 
    0.129372618974013, -0.203023536025629, 0.0407379278111141, 
    0.535536935161005, 0.592723815863746, 0.101850343978455, 
    -0.238513552406019, -0.105044778222223, -0.0422171026154608, 
    0.910348982339249, 0.371081002707003, 0.0457907941478934, 
    0.21272767402402, -0.0335166522828595, 0.0951757735402279, 
    1.1323144525495, 0.187572891875006, -0.13318128413834, 
    -0.0517537643959458, -0.0469451646352781, -0.0643800951151872, 
    -0.0520052821380185, 0.0481182102880423, 0.0523472824106337, 
    0.0240737422747069, 0.0113357781253406, 0.00404905005898609, 
    0.129350896105314, 0.0838326680048733, 0.118928832873795, 
    0.218356899661978, 0.171059608933416, 0.0286459535691125, 
    0.370212572919542, 0.391870607992577, -0.0339704814025892, 
    -0.0859628044754163, -0.071228593592937, 0.0652268996103358, 
    0.06459061551151, 0.69968301761135, 0.493565013015005, 
    -0.0353993932537262, -0.424556988571726, -0.0526505430058782, 
    0.630117533029084, 0.127295309667324, 0.010952753388641, 
    0.220533279108644, -0.233554952164221, 0.350146232227761, 
    0.361798898557871, 0.274598606080169, 0.257867469608782, 
    -0.0556273244109662, 0.543920187620961, -0.0067134975058866, 
    -0.398423798160301, -0.19003387887599, -0.140588358291707, 
    -0.220680663648969, -0.104385269527527, -0.204693848780995, 
    -0.0101979909014384, -0.260184598044348, 0.0796575680486784, 
    -0.203668164591752, 0.105104990721505, -0.0169382341825921, 
    0.0569586454829389, 0.00160571743568992, 0.0377858028837187, 
    -0.0745302281383589, 0.00994908385193073, -0.0343858438821571, 
    -0.0283876183168469, -0.0261728379337058, 0.17940952721023, 
    0.0134946103028722, 0.0293901398328053, 0.401669129000109, 
    0.178467765622478, -0.0590076480271125, 0.219327248623767, 
    0.336498742403927, -0.0197765680093623, 0.169666921688755, 
    -0.544690241730922, 0.206449989047456, 0.539077563122541, 
    -0.366835647573128, -0.458817155819119, -0.187158554355394, 
    0.711833959807604, 0.119768760927779, 0.35989769096718, 
    -0.0843293745041625, 0.36523617193126, 0.167010500491875, 
    0.00169582987135733, -0.0726496758636765, -0.0912495531407708, 
    0.291980887878582, 0.0770077261561975, -0.0161802764449006, 
    0.0779719974009693, 0.29334716269144, -0.029325697924598, 
    0.00170926883983769, 0.0596777941852183, -0.104238203428109, 
    0.0501804488768486, 0.00895241362396243, -0.0488444747607357, 
    0.0121470895395914, -0.0797251734290089, 0.073455226684416, 
    0.0627998899692017, 0.0554173300982321, 0.00936644068094451, 
    0.10783286069368, 0.117674517458239, 0.0530776479084362, 
    0.0161934696969098, 0.151931557214258, 0.155122079274816, 
    0.0493559387530016, -0.0654030801536942, 0.0589022839086371, 
    -0.0837248903251654, 0.00442914366785514, -0.0306878979560411, 
    0.0255510519410777, -0.0856870509755832, -0.0258647267408301, 
    -0.125683552734079, -0.108162036172857,
  -0.021486497977544, 0.0524678817597687, 0.0910469858139598, 
    0.0895303824482133, 0.0619976708452772, 0.0568913662849881, 
    0.0501081401234675, 0.0858306102417363, 0.115443244770646, 
    0.0988552242073862, 0.145139729738902, 0.00851322348639076, 
    0.0843444684909837, 0.431071168317957, 0.233193239097454, 
    0.0620678646977798, -0.0188494622299971, 0.282559785353719, 
    0.306549432627613, 0.211306547366658, 0.13372415273636, 
    -0.13272285626113, 0.739652095163406, 0.4683453013572, 0.440204850069099, 
    0.411908455326888, -0.0180195500985508, 0.491960940435277, 
    0.243116752780371, -0.119929080897803, -0.181067291070657, 
    -0.216285519009555, 0.129758239053094, -0.189683339796796, 
    0.0438195473472212, -0.121848878377867, 0.0170205511439617, 
    -0.0733773722496159, 0.0531392084396607, -0.216857485428367, 
    0.012333519849535, 0.088578624878917, 0.14434350155647, 0.1706774642607, 
    0.171164646143186, 0.152469104823389, 0.177430491779225, 
    0.223994801820687, 0.193493740236997, 0.121490008501543, 
    0.117266893743841, 0.133628978768995, 0.131842709713626, 
    0.170718024274085, 0.200683493929454, 0.119838413685257, 
    0.140959243129276, 0.326688731427215, 0.133001058500433, 
    0.070346358129001, 0.169907007443253, -0.260105533594162, 
    0.337391988503238, 0.43447836756343, 0.122143458948387, 
    0.043351844422828, -0.254754615651009, 0.294724255577512, 
    0.446210319110262, 0.224878450700802, 0.0355347832694565, 
    -0.225704239138138, 0.00317169147687581, 0.368821813657602, 
    0.206215946372739, 0.163853284328004, -0.0666520063275879, 
    0.451906963879049, 0.0628519510051816, -0.0656598700391469, 
    -0.395401231775531, -0.0283896296316036, -0.215141253070042, 
    -0.27693575599032, 0.15718258575099, -0.202238153230677, 
    0.0902443869907939, -0.0273668848910211, 0.131092972378853, 
    -0.230678971125242, 0.0774296371115759, 0.104985303596619, 
    0.109710724041744, 0.118015329846071, 0.139742669509607, 
    0.141627665379987, 0.140531068507562, 0.138365009172832, 
    0.152376648253138, 0.153500425389452, 0.141987151736891, 
    0.117378940053216, 0.113303899098967, 0.111620711222733, 
    0.116248473661437, 0.0985099989037825, 0.0903867309904622, 
    0.149754214614961, 0.151960749811024, 0.0755543560579631, 
    0.0368747249751082, 0.0110976040572892, 0.308065210945243, 
    0.305815741425112, 0.125099899662331, -0.0358271578056248, 
    0.204825107759651, 0.275515321627905, 0.16081815966038, 0.37476110894074, 
    0.383489173881726, 0.004612295882165, 0.452709304086057, 
    0.514768935574894, 0.311672103756231, 0.648532259628242, 
    0.48434884812203, -0.0925692587176126, 0.527277751233475, 
    0.422710154240023, -0.0382285953488361, -0.00588011577117521, 
    -0.0955660037074391, -0.147412176657864, -0.119871984029918, 
    -0.16576094663391, -0.149837696075284, -0.0455825307666635, 
    -0.0446303805529879, -0.0994876610853091, -0.108827798524284, 
    -0.0393278953346444, -0.0431372422251989, 0.0511400736909404, 
    0.0432033906924008, 0.00331566876755238, -0.298285814156107, 
    0.0609047391782014, -0.265357471845969, -0.197432299971691, 
    -0.0239884100177824, 0.0128897733763422, 0.0369750502943547, 
    -0.0254605210207973, 0.0165593815206591, -0.0125471248299974, 
    -0.010519510200456, 0.0258594051267428, 0.0489971847099133, 
    -0.0498894332973172, 0.0539399228234491, 0.0778486938279148, 
    0.254325046209697, 0.206499806738861, 0.00965939961087099, 
    0.117055933870536, 0.396408712582059, 0.133798513513866, 
    -0.111800800169012, 0.295869054980223, 0.394989473225244, 
    -0.084590615667877, 0.211098367345174, -0.536340924896267, 
    0.308948330564229, 0.587722514341883, 0.337075540733099, 
    0.195947755126826, 0.793947423072329, 0.113397292394813, 
    -0.0922127601727599, -0.123038238017984, 0.35193311752393, 
    0.130401843389178, 0.0297415707521113, -0.0147021816187822, 
    -0.0205898273064286, -0.190747567054541, 0.31607106307916, 
    0.00750019338002347, -0.266544175256812, -0.191939831561797, 
    -0.24105806409348, -0.200602515393308, -0.131806048381054, 
    -0.265583419488154, -0.0675587847723139, -0.270225598838013, 
    0.008321824492318, -0.232585293587799, 0.0477055189136787, 
    0.0718861428040394, 0.0696345464618542, 0.0602112528937636, 
    0.0837636079183271, 0.0565544245655215, 0.0914136563112251, 
    0.0622498765233338, 0.0794504660796692, 0.0921797362387631, 
    0.0193552144659782, 0.0159811804599745, -0.124968344271684, 
    0.00734708913499696, -0.0482390607413142, -0.101150682771326, 
    0.0322290350574608, 0.00239100070286347, 0.0481806472513117, 
    -0.0976824492158246, 0.0252263120316472, 0.0418130733099328, 
    0.0270573556224505, 0.0326480026780743, 0.0837536724296944, 
    0.0721198613942426, 0.107922790989606, 0.188126833145936, 
    0.0764458683950632, -0.0780571567728916, 0.38819381249897, 
    -0.115416434280303, 0.689121550676723, 0.702641357006299, 
    0.18670384537597, 0.0288064310870128, -0.140927657690007, 
    0.819839448726063, 0.573944389813662, 0.129810743518842, 
    0.000526459947393643, 0.199757227305246, 0.470451724353098, 
    0.189873079337083, -0.0858190908878652, 0.07024207365974, 
    0.529725523947241, -0.024973739341839, -0.276625564299901, 
    -0.212945353602463, -0.306266880614938, -0.23148361933849, 
    -0.206721681037932, -0.323074278260912, -0.122147823993099, 
    -0.267926131125783, -0.0801009601051941, -0.261778083793329, 
    0.00237967918318974, -0.24733898915223, -0.0363309121589797, 
    0.0577898102976587, 0.172350835279449, 0.183335702852287, 
    0.157168370531016, 0.17454165494898, 0.18665519608001, 0.150015253381957, 
    0.147984772886715, 0.198982106802468, 0.180240212132628, 
    0.142437962169805, 0.101887088983264, 0.105881000045318, 
    0.125743441241838, 0.115047858604421, 0.0833224815001618, 
    0.121301504929481, 0.108221428660154, 0.0313954080878788, 
    0.107465033809377, 0.198444752955689, 0.128188817300396, 
    0.0288522129131765, 0.193537107460276, 0.333621800930872, 
    0.163122241512601, 0.0487406200572775, 0.333350344579383, 
    0.281013073715616, 0.179390161064348, 0.0342000397831406, 
    0.645371352090235, 0.258876063721327, 0.0919237675282291, 
    0.160827526710808, 0.0559024047542115, -0.185850947433202, 
    0.768181025467136, 0.520922041720901, 0.141963625461982, 
    0.282052956564868, 0.29352427432015, 0.154181016553837, 
    0.190877342573037, 0.220939677684024, 0.258742900591656, 
    0.174549075691707, -0.0644025923095777, -0.000440447185304851, 
    -0.121338259038058, 0.114849855972432, -0.264650220332046, 
    -0.0293850901493779, -0.167218730839091, -0.187006280631639, 
    0.0382301498337782, -0.101321646633556, 0.0463695282815269, 
    -0.200995950057777, -0.0228820679681676, 0.173872030917887, 
    -0.000785162167070572, 0.230912418184618, 0.2697983624652, 
    -0.00384732129632283, 0.103231096507913, 0.371101380825258, 
    0.246813154120413, 0.258878252979561, 0.31052222468712, 
    -0.305258063319855, 0.591196676769237, 0.408193165302576, 
    0.0314888316888739, -0.228326701463837, -0.0895884208970377, 
    0.694772908359568, 0.368735548026703, 0.141739991848677, 
    0.228403892084301, 0.19258744863615, 0.00242154061640201, 
    0.0672051776544441, -0.191871333096541, -0.0320904593339461, 
    0.160119609013097, -0.100442475530061, -0.142955385989583, 
    0.0407887739636289, -0.312579734014996, -0.000679797014164929, 
    -0.327627532950854, -0.186144659351633, -0.126021683847858, 
    -0.242058476917276, -0.0969479220000893, -0.201979078901644, 
    -0.0566952378621874, -0.181030738469094,
  0.39621333630004, -0.182748380506522, 0.117982926866927, 0.640267053962599, 
    0.348958123656663, 0.416682915483674, 0.441832218829587, 
    -0.051103003720703, 0.601369460144409, 0.388657840471385, 
    0.0111147791774288, -0.16741104967184, 0.305656976117814, 
    0.0901170136716211, -0.0683490669193658, 0.133102466130549, 
    0.223889743795947, 0.0603513760264327, -0.0439808215836059, 
    0.151992016447285, 0.189346553104143, 0.110159979734983, 
    0.0703779247196976, 0.0638413224901044, 0.0886660076068154, 
    0.0750248423765117, 0.0338858761875688, 0.0447115334492935, 
    0.166751892628874, 0.154677302258476, -0.0779595839789022, 
    0.311552317624823, 0.387374923524711, 0.0680861413341813, 
    0.00551974734178645, 0.0472345052262568, -0.30391385431997, 
    0.413698944428892, 0.559012337072403, 0.116367514220036, 
    -0.033369707265592, 0.0519162746341256, 0.0243299444281225, 
    0.0328896492390772, 0.71470856143509, 0.310556416474625, 
    -0.0773280765134358, 0.395918496993398, 0.466641060267168, 
    0.0237060043775211, -0.0695181942647559, -0.0763952245843212, 
    0.00524020906269966, -0.0368102251196427, 0.0252752789087791, 
    -0.0617674571455342, 0.0496801269889013, -0.0623943553908416, 
    0.0688195308080778, -0.0382482848247824, 0.228390323499203, 
    0.0232806982406403, 0.390219308460927, 0.38461259810986, 
    0.147054773279089, -0.202887709579612, 0.491696044076719, 
    0.282730200512837, -0.220827243897895, 0.277241627776453, 
    0.632681128933208, 0.0675355832679992, -0.299506849602997, 
    0.032288593394113, 0.849927932565921, 0.175136001467417, 
    0.0756329405079352, 0.092003391193919, 0.810467974179334, 
    0.0899648647391139, -0.113529939651836, -0.0101796917525496, 
    -0.011371393535392, -0.185586200473112, -0.108295728006384, 
    -0.00666802809042545, -0.110176639680748, -0.0490653750238528, 
    0.0644902683949683, -0.191817288096954, -0.0717921501013375, 
    -0.00231194267534639, -0.0408956525969352, -0.0447388892085717, 
    -0.0277330157445111, -0.0117005904834389, -0.0385516381176125, 
    -0.0109042600131724, -0.0314527322003035, -0.0773764590103726, 
    0.0227420854351808, 0.0725498370497041, 0.0919075684696022, 
    0.0989218383146477, 0.101344745825001, 0.0770150166578126, 
    0.0985896141369469, 0.167086688896771, 0.0638585213085427, 
    -0.00588890203005723, -0.0101524845459412, -0.0408636680532133, 
    0.415064006142219, 0.417094383633323, -0.0280799348970609, 
    0.276715157602051, 0.969719437950177, 0.0698025092910383, 
    -0.114229454955033, 0.267664510083758, 0.466279341409124, 
    -0.377970735091403, -0.155960921346844, 0.935414393106822, 
    0.699821464902652, 0.346274545293318, 0.0362061763934428, 
    -0.362437849993936, -0.189595928859113, 0.53747766757858, 
    0.308868790511201, 0.19931504609314, 0.115291721379717, 
    -0.0263118677762341, 0.0900268840592541, 0.256390104184979, 
    0.310998972453971, 0.478242067222958, 0.248439420072245, 
    -0.209186096029362, 0.353395597792933, 0.411698075284551, 
    0.0664840864659511, -0.214103372130376, 0.402485421843, 
    0.514283201402585, 0.172790199886952, 0.0567478773121595, 
    -0.0944328850406102, 0.352975873821706, 0.21914406220056, 
    -0.20142429960651, 0.327280417578028, 0.556953255473902, 
    -0.088389714562001, -0.101060806612822, -0.0359248982412153, 
    -0.135565282239336, 0.727330652217006, -0.118327233240784, 
    -0.236348420494436, -0.0295475621524054, -0.457947332738062, 
    -0.168790828445794, 0.0429125025613329, -0.134940639520525, 
    0.223439751152433, -0.132948503922163, 0.0790428981166914, 
    -0.330502021499017, -0.0221176224023889, 0.0540916085843951, 
    0.107851151119953, 0.170300387212604, 0.212146514078242, 
    0.219711995467349, 0.244923454484753, 0.261667640988795, 
    0.179380023436923, 0.113089583397303, 0.396666534137926, 
    0.390932647612222, 0.169156385464424, 0.134905567807188, 
    0.431829252699802, 0.490054711611923, 0.514014515353834, 
    0.377976688802789, 0.0468755247480241, 0.0668036466930201, 
    1.01642560084538, 0.143849202499008, -0.0853188257910377, 
    -0.106652339975251, 0.441543077677458, 0.526047033844721, 
    0.406764682381472, 0.220729715026968, -0.421391011914039, 
    0.184224318382126, 0.368303355034148, 0.652816807505429, 
    0.32109552375169, -0.105847246210269, -0.0125919626009323, 
    -0.0656374855334747, -0.0639591835443511, 0.331854606504272, 
    -0.0198533166637024, -0.327483230361623, -0.228121964119686, 
    -0.0598417832680228, -0.203169651782477, -0.0741087658329764, 
    -0.182291841004592, -0.0688314214054857, -0.126446685252079, 
    -0.0404633183796878, -0.0306084840247126, -0.146165096314943, 
    -0.259936111086059, 0.139317278120276, 0.345312539610611, 
    0.104872314991806, 0.0355566596520734, -0.221165801027904, 
    0.331512894088663, 0.325889155601446, 0.130835108611594, 
    0.129917621806861, 0.457282348096369, 0.206162511822482, 
    -0.33269159545859, 0.302463125999916, 0.647226810545767, 
    0.302616642194657, 0.107096218632093, -0.230791499033001, 
    -0.0412047324899604, 0.531003940712661, 0.375130608964363, 
    0.234593836709513, 0.147627988703698, 0.101620532137959, 
    0.464074273578604, 0.46589609517062, 0.165995893382974, 
    -0.0359159365629264, 0.338210632701536, 0.489424199984504, 
    0.175162157387504, 0.0220279384893662, 0.112953565814894, 
    -0.194449338725367, 0.634694607962122, 0.315946299144995, 
    -0.0617381886843125, 0.180082185273829, 0.583024970895478, 
    0.159962025034371, -0.000725359464568642, 0.042889219672666, 
    0.0200244813478311, -0.033350585501426, 0.197418396725831, 
    0.442732200688838, 0.359851708714012, 0.0334814017152529, 
    -0.175013744522889, 0.11437661242128, -0.219795172798636, 
    0.0695219634613105, -0.358686889643036, -0.0992801344340021, 
    -0.0939141984954537, -0.216291676905362, 0.0797533853642458, 
    -0.108526561749664, 0.0973073624294874, -0.250000769973702, 
    -8.50541603650348e-05, 0.0956682466206002, 0.123705986637708, 
    0.133380708223595, 0.271321258913671, 0.338639063674186, 
    0.195628925362175, 0.0786644046559959, 0.321999534968341, 
    0.386248250889052, 0.195967866443536, 0.124008515757682, 
    0.123987081752094, 0.135075189986854, 0.144360513638612, 
    0.131002210270158, 0.141079127910609, 0.162565471719875, 
    0.159763852894965, 0.118081933021759, 0.111862889208993, 
    0.108281149820016, 0.116087126084844, 0.196740322948411, 
    0.190943262926881, 0.111152681545947, 0.0883790658168323, 
    0.211800814959319, 0.265998125736675, 0.181105653957896, 
    0.149062004835729, 0.0878351638043771, 0.284966039494618, 
    -0.285307548267668, 0.637396031174118, 0.419907710128103, 
    -0.148743969248913, -0.114345737587601, -0.157826830566418, 
    0.487282921648383, 0.0994304918730028, 0.169536725977957, 
    0.327671171277623, 0.122729036435522, 0.132760910775221, 
    0.0911912801294444, 0.0105418781132822, -0.211030040000397, 
    0.224053806560274, 0.0133731086974967, -0.126830393163424, 
    0.0750947861647584, -0.184629383793473, 0.0849199295897879, 
    -0.168445343037247, 0.111169526015319, -0.431876568665658, 
    -0.00857880165422829, -0.413106229744891, -0.285670389573982, 
    -0.0252012638865472, 0.05688953512927, 0.0855732917959742, 
    0.117202604732246, 0.174027947102886, 0.13534888952675, 
    0.118889734230604, 0.190652445119845, 0.164164352613562, 
    0.122598996819839, 0.223110566422618, 0.157920850434264, 
    0.135011483851559, 0.432062623042165, 0.336663719290529, 
    0.116621343950998, 0.219824080425554, 0.331759395710581, 
    0.234455595771228, 0.628491643837805,
  0.179447713530852, 0.115087604393998, 0.056026111394587, 0.123996159882852, 
    0.274460062872845, 0.325186429504864, 0.160420041986125, 
    -0.0388388561102868, 0.221956713627674, 0.289738443613534, 
    0.157704189438753, 0.618046633081078, 0.534213309404261, 
    0.116610733982186, 0.262376175741096, -0.060118414748329, 
    0.517251197361392, 1.03213149929035, 0.212218338381901, 
    -0.0330765209012629, -0.156810295095447, -0.102135393724833, 
    -0.118221310681619, -0.0854139538356488, -0.08598630485747, 
    -0.0485088866520742, -0.119591294764229, -0.122745118298929, 
    -0.0947998597598688, -0.0817297040932241, -0.152185207619268, 
    -0.0229403379301555, 0.0684683694177484, -0.118685748869732, 
    0.158709181458025, -0.0388369879804293, 0.0325799049129729, 
    -0.00382624893419928, 0.0462177753906396, -0.14807355599385, 
    0.0309617505830192, 0.0677529267901028, 0.0520459682126518, 
    0.155016447290406, 0.193536989336927, 0.0931929803486725, 
    0.0386446787268435, 0.262767321153592, 0.276855342093341, 
    0.133839919745431, -0.179596143075157, 0.324657392842406, 
    0.476561345209177, 0.168618178409292, -0.232885266899703, 
    0.332189586790472, 0.579612924561141, 0.257026192834796, 
    -0.156442312367158, 0.528856243914765, 0.326586669208383, 
    -0.0130725372693612, 0.530643761175656, 0.353682451541512, 
    -0.0610385115825083, 0.0987137190542801, 0.614327865746063, 
    0.166299703661095, 0.0986137897214403, 0.14766138405552, 
    0.0807690258029748, 0.267221686971273, -0.0880019172625679, 
    -0.264369315212399, 0.0664626427761669, -0.159974967390324, 
    0.196254026753998, -0.00478584267690763, 0.0922970078014855, 
    -0.296036100248031, -0.351007503244637, -0.137868281751645, 
    -0.180836767509696, -0.224265558981422, 0.122584622660148, 
    -0.270318555468301, 0.139544952392871, 0.00678460838979847, 
    0.132283250862432, -0.172894689388763, 0.0392980849791742, 
    0.19705122058366, 0.14787592949877, 0.160558621565539, 0.269158326437735, 
    0.217357032631792, 0.117404456367352, 0.108397174852893, 
    0.210346223135577, 0.301890307795672, 0.32891394762812, 
    0.268576959823778, 0.249130057408585, 0.26974346913141, 
    0.244177338542394, 0.146578197170246, 0.181290884928698, 
    0.450207538632729, 0.250706513877617, 0.0319261642810424, 
    0.250564007499335, -0.014849651125202, 0.229998445931452, 
    0.827888453099857, 0.295543633423534, 0.155436580402114, 
    0.260138765493555, 0.0952110064837007, 0.580335408908332, 
    0.249869629060265, -0.0422909482677715, -0.0204021198566775, 
    -0.00935099578560159, -0.0299980808466873, -0.00220249508033252, 
    -0.0379877391462105, -0.0160108852642046, -0.00901953735095112, 
    -0.0301282192471007, -0.00874612425595174, 0.0490695858509087, 
    0.0825483129245438, 0.0608261050537495, 0.0658416873507538, 
    0.0433870041611219, 0.0526762416021902, 0.0590527387708133, 
    0.0268317277420057, 0.0894694825734281, 0.0721839871776355, 
    -0.0272211160453002, 0.0336244242524619, 0.0824597417783307, 
    -0.044990510848512, 0.0972897885166513, -0.12446505833555, 
    -0.0769868570754487, 0.0763963650528165, 0.225604606113538, 
    -0.131062827059188, 0.12556264158647, 0.225326543442309, 
    0.157357449583897, 0.594837110341046, 0.38037721607662, 
    0.102771730258901, 0.110024210968923, 0.108393696157192, 
    -0.39190469825857, 0.148797197907891, 0.440935190246139, 
    0.121676081196234, 0.0401697223939113, 0.00168494431414525, 
    0.288471645574006, -0.0132033559727001, 0.265209972615774, 
    0.471047852955732, 0.0216581234718357, -0.0450927847816311, 
    -0.114197725486064, -0.225136519027032, 0.0877625158918678, 
    -0.176935126095529, 0.0758433988797847, -0.191151318150686, 
    0.0630738604437576, -0.163636838489133, 0.0674029819092053, 
    -0.17498541451194, 0.0699017887968098, -0.142346851196037, 
    -0.0424086228648246, -0.0839833212379876, -0.0764115159749441, 
    -0.0443157740636001, -0.0464227388276804, 0.0524296206164793, 
    -0.188095021166897, -0.102347486613298, 0.343093435947799, 
    0.136372066302686, 0.112589102060985, 0.184348015035723, 
    -0.453534338639819, 0.173728213133166, 0.684100980471821, 
    0.047531729189074, -0.0724759287916312, -0.241386155956097, 
    0.543813524536782, 0.383103318398367, 0.0946199489440396, 
    0.00887444187508191, -0.0292226736564901, 0.638349358599357, 
    0.498557165474067, 0.197172111675913, -0.0257211854773661, 
    0.756018235706886, 0.102064394576555, -0.00445922488778809, 
    -0.00998194721641214, -0.0180900262776236, 0.000467863217808409, 
    0.000536721448163788, -0.0163288325027435, 0.00685301953402161, 
    -0.020176161600982, 0.0570226864537225, 0.501172724502164, 
    0.0312648064531615, 0.0271495973070059, 0.252072750954694, 
    0.399186198220479, 0.797215726540009, 0.463405494160847, 
    0.130593403352974, 0.596212639627349, 0.319895590079189, 
    -0.00113140990652144, 0.201138658487908, 0.377692754245833, 
    0.0945268369378467, 0.263789547754041, 0.486799638873362, 
    0.130129694947792, 0.110247402480698, 0.640860792591663, 
    0.199358055662812, -0.0171375219312929, -0.00133874620788706, 
    -0.00156595012931611, -0.0033675843890003, -0.00207625069689386, 
    -0.000557612646536157, -0.00324268155539627, 4.94676990479004e-05, 
    -0.00977424870826733, -0.068413967074936, 0.301405081436967, 
    0.136086037856411, 0.0394323059724688, -0.147653297244384, 
    0.500161591549321, 0.342242353610786, -0.183936000647646, 
    0.643582766965676, 0.475176164338239, -0.130269468379488, 
    0.583481757458471, 0.422728954210805, 0.0246028143975918, 
    0.458302156855596, -0.462647836256508, 0.29456829479427, 
    0.711832408742683, 0.422117794627441, 0.0092968442282387, 
    0.562599589552399, 0.580022258165133, 0.192236451298503, 
    -0.0778942090417505, 0.242929853376843, 0.334919632364458, 
    0.152993016182115, 0.0488352070539873, 0.0208830109160709, 
    -0.234698988208903, 0.38149727913717, 0.251374942516925, 
    0.00930274536523804, -0.0684760089611799, 0.107295070976965, 
    -0.177072696927521, 0.20863419977512, 0.422564528707241, 
    0.0561014008300055, 0.0566241055296293, -0.237369137967853, 
    0.0997443569531346, 0.449415924452826, 0.139437480169169, 
    -0.178705827389422, 0.0348815629369062, 0.215077496472132, 
    0.314646215079418, 0.554211234142036, -0.0204192903548805, 
    -0.171174572641638, -0.0976710557752615, -0.133725367933618, 
    -0.0834691706138187, -0.143557639126162, -0.102857788261277, 
    -0.102872203881228, -0.105858226370265, -0.120376761054325, 
    -0.0677876297605827, -0.0961809868925155, -0.0183265014765523, 
    0.0794502854259701, 0.0486094400321661, 0.0673773036027642, 
    0.034066487601825, 0.0515964891289523, 0.0462106623580999, 
    0.052469509305443, 0.0793204577466037, 0.0229040024525461, 
    0.102796978634838, 0.107558790956103, 0.100113288554586, 
    0.257519195423153, 0.216165578829334, 0.0189698234431029, 
    0.262127359290884, 0.360218595581063, 0.0605305533014188, 
    0.082605559407626, -0.119444591339243, -0.226993652829212, 
    0.638255701615509, 0.478122863590701, 0.0489385760584862, 
    0.727360925701274, 0.404889847397019, 0.04843624234799, 
    0.710996124933727, 0.335897037907775, -0.0454319672280372, 
    -0.143495212003561, 0.500597054883679, 0.389031839749217, 
    0.308615860433733, -0.0708492170343986, 0.398645825071599, 
    1.22160220767698, 0.0492044503209737, -0.144040575339005, 
    -0.180204679263679, -0.106381197175797, -0.187408447236351, 
    -0.103113522884877, -0.167808254362041, -0.062401985453378, 
    -0.188652019376867, -0.0849124656345135, 0.0087058049099675, 
    -0.19714434672484,
  0.0384921307819831, 0.0379982970632358, 0.159284199664576, 
    0.119618210189723, 0.0310017999756635, 0.0825598147141284, 
    0.176350891263916, 0.129514306388151, 0.119790268723434, 
    -0.0584358696752115, 0.54053800730305, 0.329606895918633, 
    0.487278341854694, 0.275002094170333, -0.265922540506981, 
    -0.0409714502846105, 0.457928909221286, 0.19182257009355, 
    0.922563782247318, 0.427162879225301, -0.241384975639965, 
    -0.0847358731841777, -0.0605709813864579, -0.140898269762002, 
    -0.0444933537946015, -0.125993729932019, -0.07254201020341, 
    -0.0838597637125761, -0.0276045972635367, -0.0715758629604398, 
    -0.0655040849644557, 0.0404119838477517, -0.123928331869166, 
    0.0103471547278907, -0.0175800997617542, 0.0467487872005483, 
    -0.238981718724775, 0.00535949050637444, -0.120277650176831, 
    -0.167172184335934, -0.014740310539883, 0.0448631454331495, 
    0.0695018273461621, 0.0613424919843065, 0.0641720421509799, 
    0.0578074023931188, 0.0614364905563846, 0.085857716883186, 
    0.0746556403477011, 0.0187428385010271, 0.105455604243019, 
    0.156747854622248, 0.129002819286915, 0.152587176827387, 
    0.283514161662392, 0.232032083060461, 0.0856964557456083, 
    0.0769714625064962, 0.36036581066689, 0.23726883828454, 
    0.133265091041053, -0.171983461067031, 0.271390414990796, 
    0.502527176366809, 0.158117392294285, -0.0211269934802512, 
    -0.0698329402041299, 0.0373323328435688, 0.461347949420923, 
    0.547625829172177, 0.13435716921574, -0.220797186811027, 
    0.137597753498244, 0.370175518972869, 0.261164531579596, 
    0.174865966608513, -0.125643806261227, 0.502211204378488, 
    0.248006575210228, -0.0152008207957053, -0.264952079779102, 
    0.045610110501469, -0.310169568572786, -0.0821081430499319, 
    -0.238439324330344, -0.153456247095551, -0.172772685495603, 
    -0.182654217483936, -0.0144044659352136, -0.226553878836707, 
    0.0789940614512183, 0.00457810784511493, 0.0598962822224365, 
    0.012326411376761, 0.0566409771554688, -0.0518672158061082, 
    0.0401159997631007, -0.0177882878601186, 0.0184427204255805, 
    -0.0589382190039918, -0.0229801152137516, 0.0587399185510747, 
    0.0643628955617734, 0.0522587759384287, 0.0340411144614617, 
    0.013951806715655, 0.102231023739374, 0.179134645147685, 
    0.147056996016576, -0.25333287079756, 0.190597968033106, 0.1225695006175, 
    0.885358675162499, 0.594594578560781, 0.0653754837721345, 
    0.776918437510022, 0.363206198335634, -0.145501203672839, 
    0.488102884393542, 0.5339870203159, -0.0978927239490162, 
    -0.0769167921155413, -0.0730571657168001, -0.17691043338407, 
    0.0376534652020617, -0.133976696430454, 0.140406109504941, 
    0.0578590182842139, -0.0301331117232548, -0.0782891564909013, 
    -0.10430027281153, -0.30664964529467, 0.0145472401173719, 
    -0.122111133441124, 0.0544443310897845, -0.336896535789498, 
    0.0629229242208664, -0.197205656468055, 0.00201888537815992, 
    -0.323091952663542, -0.0496102964386844, 0.0310345679947945, 
    0.103931707655803, 0.158870651067158, 0.177444686242678, 
    0.136185299395586, 0.0849515629608717, 0.041605004300031, 
    0.127672771890909, 0.176867225066604, 0.146312002798801, 
    0.130320720563824, 0.0996902814955084, 0.103284793315138, 
    0.127640672167391, 0.112572076841879, 0.118274889274742, 
    0.134620605684799, 0.130566492952586, 0.0893673932978771, 
    0.10712149678536, 0.12119137305672, 0.114504846930827, 0.157011301513908, 
    0.183256584963164, 0.123113473905904, 0.138847960695705, 
    0.251817874403032, 0.139886081984684, -0.041893883054576, 
    0.503129414853039, 0.308573998215986, 0.085514072184096, 
    -0.0420721002160326, -0.0386942426953082, -0.0223709814594256, 
    0.707632827077864, 0.363110565278424, 0.0198381152509897, 
    0.308901118221591, 0.403303520998531, 0.162759695130768, 
    0.127104348103125, 0.217488098925238, 0.163839798761443, 
    0.546117786800879, -0.0544991436225953, -0.137229890965725, 
    -0.0353521586191067, 0.0197614157714183, -0.000315360509913307, 
    -0.266813340325165, 0.152371152152372, -0.0999358290069175, 
    0.122785765765985, -0.283129766442694, 0.011944240678391, 
    -0.156147154364114, 0.0100020197767251, -0.361949961634595, 
    -0.0357760435331089, 0.0556047683043529, 0.119215553156409, 
    0.170808497163977, 0.191951264288722, 0.156803188238849, 
    0.144848041175956, 0.204631199594138, 0.204820719775477, 
    0.163063714435378, 0.194970411708569, 0.146356641390105, 
    0.17776559014264, 0.366696552346505, 0.352494995058476, 
    0.194398221163371, 0.117486626896047, 0.244376380241373, 
    0.295700281419663, 0.362232837298991, 0.49777236191542, 
    0.312350054004297, 0.059425571301204, 0.0300543072031136, 
    0.556041686139332, 0.360941559621997, 0.145994762217242, 
    0.181563833945596, 0.129769747191199, 0.302291776476029, 
    0.675370978421722, 0.316497903496209, 0.00886469683818319, 
    -0.307170036285305, 0.0440948678192218, 0.704148919327354, 
    -0.0237061208958583, -0.178208359849976, -0.00292059735255795, 
    0.479680449917226, 0.00549689791629282, -0.158094880698052, 
    -0.00793269740815655, 0.428897061137021, 0.187725477926406, 
    0.0882042997857629, 0.0362485596617402, 0.543331690367714, 
    0.0439010564807935, -0.0180524940238191, -0.26441057643583, 
    -0.0460440566138075, -0.226850399542122, -0.0859757900558094, 
    -0.20861156130957, -0.103639843145204, -0.167823974859204, 
    -0.134064639335271, -0.0813325128608961, -0.152470362794899, 
    0.000598023686233948, 0.0623564890197218, 0.103936974417118, 
    0.0982025178602301, 0.0560373551510931, 0.0728741032200467, 
    0.0581636018323252, 0.0978459654146811, 0.125828263655623, 
    0.0588509034809335, 0.106082673275311, 0.110370901994547, 
    0.152938591197191, 0.269430267421091, 0.196970900774923, 
    0.0799448186192882, 0.235342001264019, 0.248544687469972, 
    -0.0206444958157202, 0.402828828262852, 0.410690264594714, 
    -0.0741015891373162, -0.102391403655962, -0.10237213227993, 
    0.603548273460235, 0.0161246677706881, 0.931454972562373, 
    0.653411132718333, 0.0741844302778184, 0.213229786631861, 
    -0.300557636692207, 0.105905433096409, -0.242896382156976, 
    0.0123947847973035, -0.170356846232122, 0.0313262960829999, 
    -0.241130961741798, -0.0730276540375709, -0.243928034869947, 
    -0.227321410173967, 0.0334063557355406, -0.0675807269724328, 
    -0.146387848535347, 0.0156337989611954, -0.119121077907471, 
    -0.171492042664307, 0.0904113546143818, -0.0494796799557206, 
    0.0294051258416497, -0.1542584701654, -0.0127139687343511, 
    0.0185609572205237, 0.069295305060146, 0.069856558053982, 
    0.0671790355366899, 0.056064892042642, 0.060670655093885, 
    0.0851039269655111, 0.0657400119450146, 0.0151815227578828, 
    0.100212386781281, 0.134262003819701, 0.11569949613139, 
    0.161619316909652, 0.240305379594996, 0.173575967211293, 
    0.0925933573894923, 0.137964448523258, 0.148794305486726, 
    0.145028722682501, 0.375438615420651, 0.352335077162149, 
    0.133963273947188, -0.00131930010442965, -0.295694093421053, 
    -0.00611182966805222, 0.608169803613579, 0.388251419771059, 
    0.154518516697274, 0.0562956168984996, 0.215536381298925, 
    0.144391829118562, 0.00573806925381767, -0.0130871482037714, 
    -0.0121061695167853, -0.0119375803927146, -0.0344646410404296, 
    0.0126136021506522, 0.0145208102470757, -0.021367865376262, 
    -0.0167821917777129, 0.0209574234626351, -0.0495066088209557, 
    0.00851144375476758, -0.0102539471363293, 0.0241157619079168, 
    0.00222973598282615, 0.013558043753379, -0.0915077881221136, 
    -0.0268801372132078,
  -0.00564407113790479, 0.102745341173833, 0.118898903429655, 
    0.0778790251110466, 0.100987425266501, 0.0815802947391081, 
    0.138866720324899, 0.207453836633277, 0.159823082358377, 
    0.100989445626838, 0.12039587050065, 0.133131499664947, 
    0.139319766475686, 0.152974022310957, 0.149105728350912, 
    0.135471384925794, 0.232051321123283, 0.176814296407781, 
    -0.088903295144407, -0.0108525292608237, 0.427002271245049, 
    0.505850436241466, 0.235720892086558, -0.330678733944102, 
    -0.108705658695033, 0.514164368427657, 0.252634488463849, 
    0.583768517576908, 0.763352392851573, -0.218188383152822, 
    -0.207534036839237, -0.149494614099686, 0.388733439909966, 
    0.211839761857445, 0.276473789496161, 0.33922891330246, 
    0.111749157598367, 0.565289034518848, 0.358753958865882, 
    0.0507644778902457, -0.058069038383794, 0.0873647765606342, 
    -0.16306057161608, 0.0475088184726789, -0.148159917851951, 
    -0.00716464150665029, -0.132768296144571, -0.0208964702201444, 
    -0.0778530760685157, -0.078347209117906, 0.25486673542161, 
    0.132873446695196, 0.157954629329678, -0.240510970155391, 
    0.419132644238228, 0.392971996924114, 0.14724619789046, 
    0.118578812951947, -0.130982354789772, 0.240799316704865, 
    0.877949005981342, 0.15164567455349, -0.0929620538093829, 
    0.0222769709650545, 0.0699793264842312, 0.250354858600455, 
    0.906630797194755, 0.543185803446403, 0.107994930088189, 
    -0.232239526072884, 0.324450806589173, 0.408082460146571, 
    0.0233111399002732, -0.0913180390752996, 0.0761759764643731, 
    0.180736663528048, 0.0581543316298198, 0.0248293651193954, 
    -0.130545814008304, 0.0156605655757765, 0.335133289720706, 
    0.155564147440511, 0.0626499791065436, -0.119097130276604, 
    0.0251624589710026, 0.254232965505423, 0.373143224639453, 
    0.319588505714456, 0.117747336361542, -0.170997751586322, 
    0.136310987908039, 0.377642605623602, 0.0955682579776057, 
    -0.0894702677019146, 0.194861030202337, 0.222098729526666, 
    -0.0836480074908673, 0.233006588795765, 0.391805042926449, 
    0.0581338590558372, -0.0886706621220081, -0.0262389312118048, 
    -0.356941630689365, -0.0642224889408587, -0.0556623174556119, 
    -0.24925223721343, 0.0663240920064992, -0.0699766968477911, 
    0.0432463581238887, -0.240470050774287, -0.0114981144617935, 
    0.0583410015250936, 0.0958278324331525, 0.11922236161989, 
    0.119526823385052, 0.0782470573217087, 0.0754739190397425, 
    0.113786269849427, 0.10662601630722, 0.0587896999714574, 
    0.112589251509241, 0.13321878338995, 0.134263888148199, 
    0.201344248295363, 0.216464754766514, 0.109284007950643, 
    0.134345511857246, 0.413099775294501, 0.14375857349275, 
    -0.10647089371853, -0.0296696137319741, 0.448310219392593, 
    0.329320055946668, 0.137461839589162, 0.0918181986693883, 
    -0.253221992675137, 0.423171480751042, 0.369054005998346, 
    0.160483339952809, 0.0726184790513511, 0.0962399021670643, 
    0.223704666788366, 0.107027099587135, 0.0671837263884527, 
    0.676246833358614, 0.117495097349895, -0.0672652914973781, 
    0.0170283383851766, 0.029078277133751, 0.0182685969880305, 
    -0.00811952388606994, -0.311164625585495, 0.191480460525088, 
    -0.132266275489664, 0.0405747957543834, -0.235692202628771, 
    0.005515416365048, -0.275786045983303, -0.0240537360563071, 
    -0.34422775349942, -0.0798788046855655, 0.0172285375292723, 
    0.116830995632126, 0.115753424105327, 0.111457391123618, 
    0.028402451645109, 0.0636075888457627, 0.0713916486848695, 
    -0.0291665237493836, 0.0209765029544636, 0.0855522391603444, 
    0.0831421663439351, 0.106023461993829, 0.153280882715404, 
    0.13493513345244, 0.0901471683391265, 0.0905717541133046, 
    0.148019184325824, 0.242478607207279, 0.158480041396886, 
    -0.103137203359253, 0.172633374133556, 0.440106068731008, 
    0.168930582402619, 0.0671962984526384, -0.238899636212699, 
    0.0661445745754632, 0.558738878209077, 0.196176791722017, 
    0.199270584940695, 0.457549781657987, -0.0770395194107397, 
    0.686888563300769, 0.579363197169393, 0.206006130357261, 
    0.0339710802953982, 0.776278065976585, 0.0698471108715966, 
    -0.209655367422836, 0.143144804471707, 0.426828369675351, 
    0.0704303845770379, -0.017072888087894, -0.0459057320438213, 
    0.138326060205704, -0.0474644900960575, -0.0860384830198668, 
    0.0326454887470036, -0.0525717310317441, -0.0995981467679574, 
    -0.0421408193635333, 0.0351866542930273, -0.0231352535033335, 
    0.0279208146100749, -0.0218223051867452, 0.020544573447546, 
    -0.048780882352794, 0.0250178463642837, 0.141538099942475, 
    -0.210190036859391, 0.190020982933833, 0.317392063162281, 
    0.0232997384105044, -0.11649644615505, -0.12493095896465, 
    0.286057159388302, 0.298371198474673, 0.453453680847665, 
    0.361916050017817, 0.0418793003200284, 0.226887359301818, 
    0.239631064901954, 0.622200619059703, 0.433992701564569, 
    -0.0721723456104991, -0.168172726252545, 0.0659889982048431, 
    0.192722809201477, 0.532741459738533, 0.0794871398256574, 
    -0.0295670621235059, -0.223918407439399, 0.153933424061235, 
    -0.0715437546436712, 0.127879187496726, -0.210313482731346, 
    0.12734130915178, -0.216505933944543, 0.056796171247132, 
    -0.262955432080931, 0.0301009665236874, -0.0106715496753567, 
    0.14760021011356, 0.324038325825919, 0.256961258031974, 
    0.120696623607122, -0.18543630136116, 0.344051916899185, 
    0.53633479304422, 0.0876733434954846, 0.014898582908621, 
    -0.0810270345111948, 0.86142084819745, 0.128116056759253, 
    0.0597838398419232, -0.413336408021022, 0.449229389825581, 
    0.691887357587951, 0.294193892146591, -0.119110641087872, 
    0.558993956395076, 0.426415069027648, 0.161775418527098, 
    0.123125973417671, -0.0320268726864353, 0.821413648871017, 
    0.15665137548602, 0.0735442735211663, -0.233230147828, 0.390275000558873, 
    0.366629939368975, 0.274398696943644, 0.150949947503754, 
    -0.218614690284188, 0.220229137701286, 0.241772701583152, 
    0.0185660616405014, 0.628916505079678, 0.167197346561504, 
    -0.0327217292852446, -0.165955861653782, 0.0933590350703675, 
    -0.38463934033812, -0.0644649473255038, -0.164222622860215, 
    -0.227976717479982, 0.0671980301538377, -0.171744070800526, 
    0.111048030175092, -0.242976895317558, 0.0347586700893355, 
    0.125409102259705, 0.0850793387343587, -0.00323802210475527, 
    0.244107224543483, 0.38643966341139, 0.176166344504378, 
    0.0427436831159233, -0.12140280489267, 0.434474956422214, 
    0.410613911945564, 0.133696261176889, -0.223178409990078, 
    0.30271843197281, 0.528525440201448, 0.246166117135912, 
    0.119345004963235, -0.266846768454062, 0.280709726271277, 
    0.580422793626713, 0.148301810871364, -0.151568574820774, 
    0.255305478383547, 0.466650919412152, 0.152749342173595, 
    0.0262596847149745, 0.674571363704325, 0.148528401321976, 
    -0.133666529066749, 0.229564435941262, 0.44636929951859, 
    -0.00638860202908649, 0.113497680096559, -0.285462849190013, 
    0.273988850401789, 0.410687522297419, 0.111686415853973, 
    -0.178997730772801, 0.0678506634941383, 0.408505139816689, 
    0.0343665234121939, 0.0407542531688885, -0.197422269495061, 
    0.017559514462582, 0.274854598075992, 0.164635932483852, 
    0.195608014457728, -0.200881724978491, 0.263264441801512, 
    0.127406471219499, -0.0666613198165255, 0.0312379060680878, 
    -0.170470567801507, 0.0357160700325081, -0.111950714873297, 
    0.0137649387993185, -0.400601375791714, -0.0841819604222449, 
    -0.196697881856918, -0.327438445197458,
  -0.258631419248274, 0.00356325250948854, -0.210237612302706, 
    -0.0895898875037878, -0.176870046101708, -0.0996337428927957, 
    -0.171354154735852, -0.0939382593082894, -0.131676142827994, 
    -0.10569321857945, 0.000326926313610518, 0.0999093249766647, 
    -0.0326908981191077, 0.0499463291622631, 0.0119952727379465, 
    0.0398931644153434, -0.0574948856427175, 0.0153867388604496, 
    -0.0241589522666159, -0.0692754229616139, 0.0407890809065556, 
    0.105302387837764, 0.075217346189074, 0.0939740581044736, 
    0.150793678330275, 0.104554129497622, 0.122945737867817, 
    0.337213079827647, 0.0886685693789819, -0.222510439976264, 
    -0.11179741817948, 0.353482040578257, 0.394035233905238, 
    0.472364090060065, 0.350360867497501, -0.0341356798925426, 
    0.425764299854051, 0.479976406684989, 0.0278744633639878, 
    -0.131956894060687, 0.671725135275175, 0.524278380606633, 
    0.167814900363907, 0.151276931333972, 0.483345631075123, 
    0.261218674747419, 0.204262002944455, 0.300107196887368, 
    -0.203165242586385, 0.0292033806465214, -0.232125411711584, 
    0.220709994244545, -0.454974523951951, -0.0602784861958519, 
    -0.258980212726273, -0.282204718134731, 0.0518881833858498, 
    -0.318238317781898, 0.0794633404063649, -0.283204524903397, 
    0.0279676343128574, -0.0199452928116808, 0.0437635350924385, 
    0.0267226796606824, 0.0821858374682772, -0.0270655052499827, 
    0.0530945016983359, -0.0308098351297698, 0.0090760586900383, 
    -0.12563152508266, -0.0451677355988837, 0.0454392874303171, 
    0.0465127761597944, 0.0215516752469286, -0.00921815851357585, 
    0.246830319637413, 0.05283922255336, -0.141818243706197, 
    0.0627092990949111, 0.18794006347314, 0.146912331071008, 
    -0.218554640401983, -0.0298352442910106, 0.971019509388106, 
    0.281354198127947, -0.35730486182706, 0.185357251312124, 
    0.634708742355835, 0.326053610603335, 0.203550086931411, 
    -0.132982758849065, 0.557752004424124, 0.219134600908571, 
    -0.0024152011353273, 0.034968508915317, -0.0448918157487883, 
    0.375026753366041, 0.867909611398265, 0.0678340463664744, 
    -0.110569685635434, -0.0605042618359848, -0.293145730966493, 
    -0.0335075660857574, -0.248039934912654, -0.0654051886409865, 
    -0.289845312679039, -0.029793751546616, -0.239053203316831, 
    -0.0352713168072328, -0.231683230536107, 0.108979301970125, 
    -0.006374326511618, 0.0514683861194684, -0.0112734522205786, 
    0.0149879890982876, 0.0185931241369173, 0.0234211874067874, 
    0.0726362074447792, -0.0130531575872449, 0.0663969022673718, 
    -0.0981891706379191, -0.0246094895242025, -0.0272635586503471, 
    -0.0458753366897814, 0.0131701092941481, -0.0424880344889562, 
    0.0169982353125837, -0.0125433291367052, 0.0530496852530834, 
    -0.0901138806871413, 0.0292977561795735, 0.111105485137362, 
    0.0906991669132517, 0.0649930571187983, 0.0102372554583485, 
    0.298138897548896, 0.172701541839928, 0.0379161220324836, 
    0.123433397767227, 0.0566355647735801, 0.0955686634174663, 
    0.574983829879262, 0.289505042703467, -0.0166674991081652, 
    0.151825497595274, -0.577815188375265, 0.82162139283283, 
    0.580666048262852, 0.281889657146811, 0.453591513369665, 
    0.200664576559439, 0.000507027450969019, 0.0252580880831551, 
    -0.117310392963446, -0.016173285119503, 0.13612175227118, 
    0.137813353038891, -0.0370598194401448, -0.132110103437858, 
    0.0948403857441984, -0.351898259124958, -0.0424994408295971, 
    -0.224918904255904, -0.235766277300736, 0.12199825559584, 
    -0.184741779757854, 0.129218207651081, -0.0738962165066717, 
    0.125936262356272, -0.206701005344465, 0.0574814066194263, 
    0.0339352386171081, 0.0495005481097084, -0.0312788312926264, 
    0.0279188691118869, -0.0144801611037169, 0.0145961377540169, 
    0.0217653010202114, 0.0618295455508279, -0.0341651590958088, 
    0.0541300605496863, 0.128001121469608, 0.205213779996556, 
    0.132956678611737, 0.0218775491792118, 0.0121364298563578, 
    0.203141029512397, 0.183827483102965, 0.0457461492176994, 
    0.0739623276234866, 0.41525647058839, -0.0234215036212265, 
    0.141225897989973, 0.247331897291537, 1.44169095986966, 
    0.0191515953160704, -0.438047931187361, -0.0348878497811556, 
    0.937134858293343, -0.0396998264143705, -0.113451324234383, 
    0.0422137984233895, -0.0611232405162723, -0.0662283684223688, 
    0.0470371124618687, 0.017149383135608, 0.121726851123682, 
    0.192757876384788, -0.122114892970096, -0.0550742426832543, 
    -0.150254609326213, 0.0540852544172904, -0.234999029312597, 
    -0.0402390135898706, -0.153296899739094, -0.140163274535004, 
    -0.0222322668164157, -0.145177981425863, 0.0354221483287258, 
    -0.149913490608487, -0.00352276495274249, 0.0469571438410191, 
    0.0536239794343864, 0.0665201354609131, 0.104176946193809, 
    0.0858123874408171, 0.0478233998628296, -0.0592952885685329, 
    0.284942861907529, 0.197086420659035, -0.14015838493847, 
    0.103650312766136, 0.624350118325228, 0.135401329514293, 
    -0.0480848299136958, 0.263044059552285, 0.288201806824578, 
    -0.171038560985311, 0.953415900546481, 0.398336003276351, 
    -0.127971100777691, -0.228848072769432, -0.118135454413196, 
    -0.096151833276784, 0.838247264246061, 0.355774676485467, 
    0.00943675951689686, 0.644588385609826, -0.0878995487310076, 
    -0.360556079777471, -0.142536851146595, -0.143328259721152, 
    -0.154240994310907, -0.166175349037165, -0.120460773073387, 
    -0.151550749865814, -0.099158650395601, -0.173125803411783, 
    -0.0662031749569645, -0.112422025228271, 0.00517605871640604, 
    0.0072045766677792, 0.235793945686276, 0.243758441295724, 
    0.221038474908547, 0.239893203119057, 0.132840026405086, 
    0.0780191473710731, 0.383276358279808, 0.337924450351705, 
    0.134395270673291, 0.0926433495335172, 0.0818106141667851, 
    0.09725232765672, 0.0660732297857917, 0.084498140177575, 
    0.0797617885590311, 0.0809461145037191, 0.0347564494269648, 
    0.044686628571074, 0.060351040154013, 0.0740450901474888, 
    0.0988346739508216, 0.117901216241585, 0.12648556078502, 
    0.113757546845249, 0.0830805086624399, 0.0949791764022488, 
    0.110208145462286, 0.074200905987024, 0.122103939712451, 
    0.130319647636058, 0.173943741364323, 0.243982718585968, 
    0.185536319353216, 0.0796507827211804, 0.188400539354645, 
    0.369365067043464, 0.248622516995591, 0.0640963906999824, 
    -0.0349048972274255, -0.039044293703013, 0.61470176204827, 
    0.14283398630707, 0.141579322471234, -0.264287159881364, 
    0.164297916116678, 0.458769452787596, 0.247779667912304, 
    0.102680978881634, 0.153358441855158, 0.208961965587474, 
    0.199289481414857, 0.109825375001236, 0.244897916307153, 
    0.364542192005087, 0.0533098853082669, -0.00621581449757086, 
    0.0153416376170712, -0.074196297311355, 0.0395754062556858, 
    -0.363536393025993, 0.107896716998381, -0.0931859107144437, 
    0.0168167929630015, -0.26035922025494, -0.0271747359830275, 
    -0.112403917926088, 0.033523905791874, -0.281577367338375, 
    -0.0360134392350673, 0.121651815173157, 0.108334897438567, 
    0.146249401552828, 0.2259776450376, 0.18310503176458, 0.140312252491637, 
    0.198381751770172, 0.204091506710914, 0.183892693503289, 
    0.25881337881138, 0.198875570114985, 0.17448634903673, 0.409153795312493, 
    0.36754777261805, 0.140297339758198, 0.00523391210146701, 
    0.29194712756726, 0.63744198163791, 0.280892941011486, 
    -0.128109922491559, 0.331501651021061, 0.321164998426604, 
    0.194098306398808, 0.592987602225985, 0.225459548870641, 
    0.0129794773448257, -0.362510001621304, 0.236425154730839, 
    0.18854195916473,
  0.00529871890275156, 0.051391907249963, 0.0531592972276007, 
    0.0625130795188122, 0.00164199165530347, 0.0540797790921693, 
    0.00404470043815579, 0.0176302307352774, 0.0340233153738923, 
    0.0153053965247162, 0.27243665624793, 0.0825454759561104, 
    0.0275774665231471, 0.416441210871753, 0.244774189174327, 
    0.0821812766149097, -0.0440590874829593, 0.105701207355085, 
    0.431011433605145, 0.308733602565329, -0.0637637298761859, 
    0.82528814796996, 0.324182470353251, -0.0191261789058077, 
    -0.0225472680169478, 0.156820632507282, -0.109255086425225, 
    1.3821417186523, 0.386571679687343, -0.0533250653105361, 
    -0.125846655769532, -0.157752599146868, -0.0902674294844982, 
    -0.0797157463029249, -0.096043769640382, -0.0695833808696019, 
    -0.151671618295982, -0.0718618210167374, -0.0497800819874205, 
    -0.187185658305985, 0.0670179636205925, 0.0487148014869837, 
    0.0814199386157259, 0.0500035301422849, 0.0774203176447552, 
    0.0560047093703459, 0.0311720354701194, 0.063384101847614, 
    0.0923999206080059, 0.0926131847031527, 0.0027699133774995, 
    0.0415150604734087, 0.0280338342942225, 0.0147060043449747, 
    0.0735875216261362, 0.0192007709039488, 0.034674094627299, 
    0.0582673882232622, 0.0603289276413327, -0.000145528520404822, 
    0.0649964107935688, 0.0981930029221156, 0.112807645272685, 
    0.150875035694167, 0.170116332268328, 0.161062450178092, 
    0.196416139780156, 0.187690936531957, 0.0870425301938447, 
    -0.0711913452768948, 0.463796965788312, 0.294870743611915, 
    0.0942041565189532, 0.230289759907926, 0.0901664835750518, 
    0.227385267049459, 0.782969509260573, 0.217931125794756, 
    0.00985458517866653, -0.0718179650614878, 0.567030860224166, 
    0.202284693457722, 0.114964083817659, 0.134749440819761, 
    0.0859310614196034, 0.199633810076358, 0.206519687559977, 
    0.159495715955489, 0.926041239574701, 0.043175336277709, 
    -0.27525498433349, -0.139577637917169, -0.115521537517391, 
    -0.177103523136943, -0.128263721925476, -0.182420625707835, 
    -0.166819029542367, -0.112603360797375, -0.0585915954750598, 
    -0.191788238587203, 0.0787059593855851, 0.0146448920398632, 
    0.0628585608329565, 0.0287852850718531, 0.0569411951685126, 
    0.0171079761170445, 0.0516638212856105, 0.0458564044990309, 
    0.0822016229773229, 0.00336750118781984, 0.213892906116145, 
    0.166816608577742, 0.0669236150189307, 0.0669340627437048, 
    0.248223754827444, 0.21410318276629, 0.174338565300048, 
    0.395714813308651, 0.203798070032232, -0.0224831076186589, 
    -0.232627711676481, 0.357286026013593, 0.623623640196749, 
    0.0903242372561407, -0.22481642581212, 0.892076324926858, 
    0.666608084198341, 0.755814920564364, 0.838876126765675, 
    0.032192021371078, -0.223396723780285, -0.0396249334688529, 
    -0.124115864142797, -0.104491267355532, -0.0785793036931779, 
    -0.0751210670370749, -0.0700684166333554, -0.104725824952488, 
    -0.162587187624891, -0.023894880614078, 0.0175564285319881, 
    0.0922702499824641, -0.0229370488702147, 0.0567812754406064, 
    -0.0392841229703988, 0.00666761383445443, 0.0153512332679239, 
    -0.0109703477709339, 0.058252702970382, 0.0212281971466278, 
    0.0438974259444479, -0.0408405659340343, 0.0316821164734388, 
    -0.0165271813060407, 0.0319873565436871, -0.0449243775626469, 
    0.0218725432657124, -0.0272014794835979, 0.0196638729129889, 
    -0.062524026103681, 0.0383153660167864, 0.0404191824764215, 
    0.0923671498541557, 0.188049117714881, 0.17035162011879, 
    0.085877375347384, 0.0164333093874594, 0.18891247240333, 
    0.286838468784219, 0.129102475555322, -0.279491675270603, 
    0.28887893833436, 0.660607949615582, -0.0417952938215566, 
    0.126257126639688, -0.268420443068837, -0.0424697578152572, 
    0.708101959323581, 0.108950192270588, -0.125375064360374, 
    -0.132548412451142, -0.0732813059680428, 0.562827795227999, 
    0.371276998630111, -0.0428735575489855, 0.281020746988148, 
    0.65616137506539, 0.672585160811693, -0.0324911400934593, 
    -0.31699746230639, -0.427731254998938, 0.065390882152425, 
    -0.326504325820283, -0.194797388148042, -0.147927700885973, 
    -0.24299364008035, -0.0599563726216691, -0.234661258810825, 
    0.00794689410152574, -0.238824445755519, 0.00669328061779524, 
    0.0582455753939826, 0.0935875067630045, 0.218393187290266, 
    0.236710199640917, 0.128599903754894, 0.0662677404552878, 
    0.249231306210137, 0.265224904115373, 0.161046184727639, 
    0.122450512555343, -0.126647433813285, -0.0295080721649582, 
    0.658922096714739, 0.228834475507646, -0.0788349520981153, 
    0.241629679259704, 0.382211606191875, 0.0712098783018648, 
    0.610153110978652, 0.477501618801824, 0.0361664981771259, 
    0.00716808651384183, -0.174774229786768, 0.060495392480919, 
    0.44059121334546, 0.305211547960008, 0.650667736047494, 
    0.525577483303728, -0.0816858520450172, -0.180862482081441, 
    -0.0886361807890739, -0.184809869655105, -0.173551890452616, 
    -0.162331242233191, -0.0706424095238158, -0.191004856866089, 
    -0.102955662567231, -0.166803291856989, -0.126968009769335, 
    -0.0390758075725585, -0.00790586181446859, 0.0133221393737478, 
    -0.0444790722189239, 0.0735209947777133, 0.000521916354702806, 
    0.0505725036882798, 0.0364677188412158, 0.061773191411275, 
    -0.0540744065089718, -0.0143055880247604, 0.173494663614114, 
    0.141749208396254, 0.0115765500046615, 0.242201606240024, 
    0.184144280421968, 0.00954100258675918, -0.0127521788073301, 
    -0.0834454224779776, -0.022464497413081, 0.647515489240412, 
    0.165167348838809, 0.836331692374049, 0.802722897009372, 
    0.330046221667033, 0.261484730476608, 0.127293130373819, 
    -0.19778865120721, 0.800853765195509, 0.100087548817403, 
    -0.223643422760027, -0.123937797627413, -0.11536233760785, 
    -0.21170264003515, -0.123611586240103, -0.207453610893564, 
    -0.0666562301088136, -0.177552185121809, -0.193791535088932, 
    -0.121408154404256, -0.237498208654048, -0.0508133622245518, 
    -0.337940132315442, -0.0857179196481676, -0.155830362325039, 
    -0.255038515466242, -0.0193597036861305, -0.103457115632943, 
    -0.0607782577081932, -0.255344523067158, -0.0962921601888908, 
    0.00554391890939249, -0.0629691157411189, -0.0216413291596805, 
    -0.0239576520003682, -0.0232610380640376, 0.0781328828993755, 
    0.0217139123236278, -0.269653199329716, -0.0750744460853496, 
    0.480146488882825, 0.165459190819864, 0.689150885437347, 
    0.574647179568287, 0.0431445774265149, -0.437165187589588, 
    -0.0258237736449529, 0.623309364727534, 0.457574795906391, 
    0.193589741481063, -0.115590583017731, 0.263721477473529, 
    0.31577023201512, 0.0970711821950512, 0.0421607542413524, 
    -0.117449683319487, 0.0818758165329203, 0.25299168286421, 
    0.0507111432162342, 0.0649109963018485, -0.175442099865093, 
    0.0357784437733796, -0.273270076274772, -0.123401112689711, 
    -0.0338335463039877, -0.165861601664818, 0.039881435627453, 
    -0.148119733816322, 0.0235609451403895, -0.176300186284588, 
    -0.00451871542905398, 0.00272617651683418, 0.123099786643855, 
    0.225413911514567, 0.123193367048563, 0.010942849532486, 
    0.0701297723550223, 0.2363240700165, -0.0148975381502852, 
    0.00526519072256261, 0.583339162890458, 0.431939865646001, 
    0.289004252662874, -0.102542135885441, 0.991036780960143, 
    0.251917871288332, -0.0759676089899643, 0.491133787412478, 
    0.410506434506401, 0.0308024261979341, -0.0722204885185501, 
    -0.132437389934866, -0.0714390038543499, -0.0141640842298554, 
    -0.116126025230206, -0.0627820702711195, -0.0661715017056866, 
    -0.0233728697933786, -0.0366652024695844, -0.0435315846864421,
  0.196320420427458, -0.248602566790856, 0.291849002950161, 
    0.751016790854844, 0.238299153605833, -0.186957138331276, 
    0.505518216893693, 0.685018435906324, 0.182123736291362, 
    -0.00387070171510131, -0.101401813266036, 0.302866274906983, 
    0.705566044433944, 0.227978726032887, -0.171249335555878, 
    0.201319037604574, 0.504820837881229, 0.18479799083315, 
    0.0737007662526019, 0.154062153027051, 0.0350809835498949, 
    0.248776520438252, 0.186921228856267, 0.628413244100428, 
    0.489095425564377, -0.0823221007662582, -0.2132251373189, 
    0.146509639201233, 0.214722141882401, 0.0138703246427516, 
    -0.101946061271779, 0.25711797987979, -0.0897140461745923, 
    0.204501129427668, -0.211659034176897, 0.0803871461588116, 
    -0.153122228791096, 0.00852691271562908, -0.332621188467028, 
    -0.177901084526512, 0.0115709984819925, 0.13690831971387, 
    0.10634545308468, 0.0904315154778154, 0.0904083814424242, 
    0.109928856158094, 0.141213603338625, 0.142159313153009, 
    0.170328590311029, 0.168432184078422, 0.136219093627399, 
    0.106106040684067, 0.103212587341461, 0.105482050060239, 
    0.110654756956145, 0.0910195563333106, 0.0900446255152525, 
    0.122772648437919, 0.117196718658708, 0.0675228132488739, 
    0.108235602255014, 0.157597144145245, 0.168304627063406, 
    0.113576868968576, 0.0937652522392045, 0.274267302290874, 
    0.213745460654626, 0.0762663223561584, 0.0381221923593798, 
    0.0164851029245727, 0.636231506893314, 0.0863363958852391, 
    -0.113957168651327, 0.531863826399161, -0.161032948334876, 
    -0.249696988375131, -0.068081961515995, 0.219553691894624, 
    0.651405311907571, -0.0712193001207536, -0.201882817390589, 
    0.114778218333719, -0.0454724049828295, -0.00814101000095018, 
    -0.102350420171142, -0.112651191549472, 0.0967963832168496, 
    -0.011705515265852, 0.0107612779962121, 0.0129082625805476, 
    -0.0897882755512033, 0.0403417911688862, -0.142084982453794, 
    0.0848377488602766, -0.353960675766278, -0.0495549243021402, 
    -0.124585039570309, -0.153461850454024, -0.0674183305364112, 
    -0.183279241688033, -0.00269406544984581, -0.00857755562047105, 
    -0.00778493351710494, 0.303514806003237, 0.173868271726184, 
    0.047201277284405, 0.104132454776072, 0.254329252329334, 
    -0.129453642150044, -0.063982179530719, 0.693115389522242, 
    0.20131342430029, -0.185705561681799, 0.401079993812164, 
    0.469637698128182, 0.0661791187452054, 0.377715922768891, 
    0.721533967363167, 0.251868564846176, 0.0131249321127084, 
    0.0821358031334116, 0.455789126002052, 0.383867043255099, 
    0.238943399071538, 0.169513399995936, 0.117023331322285, 
    0.136106590088993, 0.252136127577884, 0.140862969092998, 
    -0.0620244596497731, 0.101544440238104, 0.381400418000494, 
    0.160557879566862, -0.0879014271922348, 0.256441594134788, 
    0.332800449792535, 0.101681058988139, -0.0093790111531358, 
    -0.0507271814771915, 0.251076827705668, 0.543398350567828, 
    0.277364849601123, -0.0430824398508262, 0.501375159162046, 
    0.315220724172045, 0.0904523843046273, -0.119617947433683, 
    0.432547033827323, 0.444650043244545, 0.212119515581974, 
    -0.00256412647740449, -0.000937643202201716, -0.182486636809917, 
    -0.113457863528382, -0.0548942905057777, -0.13795189242856, 
    -0.126271557643751, -0.18487739309309, -0.177086032124451, 
    -0.11109862324072, -0.0876332686347172, -0.147806499962279, 
    -0.0485252207760006, -0.0051613264375326, 0.0618296945529471, 
    -0.0961223275400539, 0.0673421255528555, -0.0874454564124527, 
    0.0327927845078983, -0.181686522145137, -0.0428538418054737, 
    0.059629500623833, 0.0641171583050632, 0.0630806406359804, 
    0.100087177724081, 0.0840060051772178, 0.119049246332889, 
    0.294140049093408, 0.123215445059928, -0.270663653206081, 
    0.0558580412661973, 0.53925273058073, 0.187457508813966, 
    -0.00574447420493648, 0.2294803514636, 0.010548917720115, 
    0.220022674446929, 0.869163328061544, 0.222450658288526, 
    0.0677874597261846, -0.263113728885811, 0.471699557922717, 
    0.336381824059397, 0.0686476914615729, -0.0293071019589816, 
    -0.0788848637733465, -0.337171025827571, 0.455855009356522, 
    0.293837386441987, -0.34150764134993, -0.367780812712121, 
    -0.255809296022136, -0.142948915593889, -0.225153816008053, 
    -0.078966944761538, -0.223766297533929, 0.0351705710429827, 
    -0.29147826057995, -0.00766467891606523, -0.202428931470518, 
    0.0336588864326704, -0.0254482972773454, 0.115374137012225, 
    -0.0688604520963256, 0.0949144546309834, -0.054951844829434, 
    0.0993220877762951, -0.0670865191923396, 0.0574705718606105, 
    -0.272682784251634, -0.0608623721673977, -0.0259068651946405, 
    -0.0236878026578585, -0.0125288387101938, 0.00890660473378926, 
    0.0196198626211059, -0.0901816462286691, 0.173315659507125, 
    0.133655413967038, -0.251571054579061, -0.107926125446572, 
    0.545739021613423, 0.134793696307953, 0.00446676376803766, 
    -0.108834483024073, 0.207295876903207, 0.0642633035013787, 
    0.546638299904223, 0.690233746254166, 0.0978939379494785, 
    -0.0323944292208202, -0.122101793987424, -0.317276123500183, 
    0.85647912780768, 0.0843595306400901, 0.0315552859359451, 
    -0.531683719465818, 0.215931352263625, 0.776496231490143, 
    0.4634563700473, 0.284832458255432, 0.367642871042636, 0.175287249196569, 
    0.0354596094296598, 0.112381206794229, 0.267030319348478, 
    0.128291300659295, 0.011373481723013, 0.330862748049459, 
    0.227908576467089, -0.100762862402314, 0.3377876448061, 
    0.407454304840479, 0.284040453761833, 0.250006834856681, 
    -0.146011566257127, 0.162939501225139, 0.312977106746536, 
    0.677034119800474, 0.246821212056987, -0.188218514193635, 
    0.104263304277676, 0.510906550660644, 0.0791399853983734, 
    0.127239947732589, -0.329370309712002, 0.46552667707645, 
    0.396898123360412, 0.226820928792208, 0.337947147343972, 
    0.133330769580085, -0.0670644789570939, -0.0905939307866997, 
    -0.0904147037610822, -0.114109466326083, -0.122079951647478, 
    -0.0972621310540755, -0.0901883778061512, -0.0420736667561911, 
    -0.188703888222632, -0.0357598034734461, 0.132735064705121, 
    0.184169271522511, 0.151240654199708, 0.122577378384371, 
    0.114224409602169, 0.0743812675702994, 0.144234169949767, 
    0.223677018463002, 0.139426506443473, 0.0685380483864929, 
    0.0728744109465912, 0.0806161472584729, 0.0751041725737948, 
    0.0845090384462547, 0.0704390847828527, 0.0724234279071631, 
    0.0860741451252332, 0.0941069418804859, 0.0539135149024369, 
    0.0870083178925391, 0.108336098367145, 0.126782329500716, 
    0.170090284154501, 0.171803904468564, 0.106012752049434, 
    0.104712452735535, 0.243347195146973, 0.160342233882396, 
    0.0517363528700017, 0.212675498623792, 0.233353075979659, 
    0.00919034885071672, -0.0379229359399316, 0.351141197402956, 
    0.389067349559924, 0.452193544304414, 0.404959129992179, 
    0.096919311635818, -0.36106492639152, 0.198008871399638, 
    0.634073725990605, 0.115425265209777, -0.114623933914996, 
    0.0986668841411304, 0.352807778605516, 0.0945905709870463, 
    0.468044030661631, 0.564355324212907, 0.0101459380313769, 
    -0.0856507770338695, -0.132535673075636, 0.0577490244522842, 
    -0.0651915844127333, 0.00637254667457275, -0.168753711883225, 
    -0.0204461398307203, -0.0777778939250232, -0.0555916428024895, 
    -0.080277340512731, -0.162081680730661, 0.109264834014343, 
    0.332328327727744, 0.133701302475612, 0.0219466019575653, 
    -0.141185761187704, 0.0722145567756824, 0.432205455794055, 
    0.409441491784625, 0.306393875637986,
  -0.0729405432941603, -0.141711856776089, 0.0259410882445248, 
    -0.0463781780931887, 0.0697550509427531, -0.115681113154182, 
    0.0739644974189333, -0.0667987096455707, 0.0379973945509246, 
    -0.160032884082426, -0.104064063601567, 0.205076254244852, 
    0.147662133869833, 0.0591602078183818, 0.0940601441396671, 
    -0.059237662385531, 0.101346006336571, 0.491461301475801, 
    0.106376283896021, 0.0552446224551259, 0.378910155326329, 
    0.158160087787741, 1.02778331965838, 0.291097202646812, 
    -0.045644650920048, 0.730125166824492, 0.345496739425249, 
    -0.102233550527193, -0.194440805698992, 0.360293023881943, 
    0.142036797607851, -0.410079977075316, -0.211205552987534, 
    0.098394206835271, -0.231450911011529, 0.0343431919513801, 
    0.0583701148755509, -0.00263997109151182, -0.123354413854539, 
    -0.188022796585416, 0.0653598763695341, -0.24576118395511, 
    0.049061552504482, -0.270624322629119, -0.0268708167637244, 
    -0.200765324163873, -0.0236635534119354, -0.168372788281119, 
    0.0121867038178984, -0.178553250956967, -0.0268191123261204, 
    0.0182710722755931, 0.0105221487294477, 0.0197702319985878, 
    0.0155278136455223, 0.0220779656928931, -0.00453366410949801, 
    0.0592332743151415, 0.0645979045789527, 0.153179550297423, 
    -0.200167243780121, 0.387595621097381, 0.390119931293675, 
    0.132872525266818, -0.0998090374115421, 0.141337424713463, 
    0.637125396498742, -0.0296517218338197, -0.114639375808951, 
    -0.201574506107667, -0.344916833367531, -0.158256218788271, 
    1.02852812383372, 0.300187412049783, 0.172699209327239, 
    0.386782206590589, -0.594363035584984, 0.433849301404799, 
    0.856367119182258, -0.335898698220497, -0.163038269258421, 
    -0.203056014627039, 0.00674646858628881, 0.101743940880895, 
    0.00190112856981553, 0.0315670889566139, -0.0156783233176675, 
    0.113618265629906, 0.0793551563952075, -0.138651726848575, 
    0.330312882586573, 0.226403813797143, 0.0896077756114937, 
    0.0633221154115682, 0.059052398252712, 0.0326621204137835, 
    0.377775041643326, 0.334782851145175, 0.17108092107621, 
    0.270232895965414, 0.326232942715678, 0.232579880179897, 
    0.137384209184077, 0.117762474920281, 0.163957289982787, 
    0.0722808740478594, -0.0651332970388615, 0.121718394317232, 
    0.241099124497888, 0.0471330762828484, -0.0519972581716995, 
    0.0228943955621928, -0.0182434240319121, 0.0287919647505511, 
    -0.129512417703137, 0.0159418753605762, -0.090123775278672, 
    -0.054569836485376, -0.0441928624947553, 0.00866190605020831, 
    -0.0264507084682292, 0.00856361425079333, 0.22199235727672, 
    0.21987459955021, 0.132204395368731, 0.0239133900872556, 
    -0.205906305302105, 0.133714369105099, 0.543352171427348, 
    0.141732841832484, 0.0186857740707792, 0.248615165403992, 
    -0.301584667421703, 0.666751738368515, 0.669959746635944, 
    0.343491988578613, 0.331052827838631, -0.26875617584915, 
    0.737787130046895, 0.826816971734775, 0.0152409327879462, 
    -0.0290190583075881, 0.112403050943594, -0.0543687432914127, 
    0.215667328118543, 0.118703228407054, 0.0645570578235594, 
    -0.121277436706712, 0.0894571309676051, 0.118407526716458, 
    -0.0227476635531028, -0.0102946114884227, -0.0264865565727868, 
    0.0388428969901141, -0.0644030114172979, -0.044070301695519, 
    -0.0687083237901927, -0.0223035695076613, -0.0892346831753489, 
    -0.0836545760272018, 0.0272536050009944, 0.0259573070887287, 
    0.0279846450599542, 0.0227178049759885, 0.0388045922936908, 
    0.0174962337559099, 0.0335652255948278, 0.0265054860573648, 
    0.0374173560896209, 0.0109541325526931, 0.0708339946871661, 
    0.0919007462853022, 0.0985203411828389, 0.117421783200319, 
    0.155650725654411, 0.123427682240936, 0.0599712388600839, 
    0.137631676400889, 0.180386770521997, 0.0898915551317486, 
    0.0954833180586818, 0.0448492374767799, -0.127248675363438, 
    0.285498803470779, 0.603157209101539, 0.147458994898341, 
    -0.0288588159113234, -0.0260680596475341, -0.251079388729058, 
    0.626607469547488, 0.380225928948874, -0.00759566637210624, 
    -0.0993025316315226, -0.0145331240242459, 1.09611934540672, 
    -0.0157711110228935, -0.553060130241846, 0.436269310023177, 
    0.524325488962514, -0.401051250514165, -0.125362236189257, 
    -0.237268438610939, -0.118693891267684, -0.318109083614704, 
    -0.140798405200048, -0.237814868344531, -0.243649358853985, 
    -0.159787604477124, -0.280427002389817, -0.109259540742319, 
    -0.0260301810255765, 0.0877504707293768, -0.0380840811674488, 
    0.0403671030569632, -0.00544146901018727, -0.00713539144542599, 
    0.0794923846170129, 0.0129936408568183, 0.0938673438784848, 
    -0.00738610944312693, 0.107474491938264, 0.0804589022001115, 
    0.0152658561764677, 0.170934298808979, 0.175234488979294, 
    0.149827907229654, 0.342158428516161, 0.130305784132665, 
    -0.0464648937911196, -0.14064847118528, 0.1688076064253, 
    0.360343507165784, 0.0339115943321979, 0.685834935049652, 
    0.341863479234427, 0.0855764969057557, 0.13473821505669, 
    0.158764208655313, 0.59589731801412, -0.0482387781741665, 
    -0.099235872164046, -0.140943498763874, 0.0183735438918501, 
    -0.0476772785970142, -0.10779335801494, -0.0706953907545173, 
    -0.124356376575482, -0.0539523415595126, -0.0783640543963081, 
    -0.0770737540300694, -0.030183972354951, 0.0279414896697132, 
    -0.119276237976888, -0.032251726594248, 0.0599827401538574, 
    -0.0580938657848572, 0.0744500170727642, -0.0152041131713619, 
    0.0250822239382882, -0.101452023272187, -0.029655215994518, 
    -0.0791264202285616, -0.0625106115930945, -0.0675448429643333, 
    -0.0445961427100446, -0.0725985068577487, -0.0515105545893572, 
    0.0584388143157691, -0.0884352228933996, 0.248470207610804, 
    0.064119335536462, -0.0279883281658277, -0.253277966563641, 
    -0.194830233154896, -0.0590893375577458, 0.974678476341073, 
    0.344567303097101, -0.0663429214121825, 0.148137400629011, 
    0.303709535177779, 0.442936662227346, 0.765280832952504, 
    0.276775428913687, -0.0929595639020754, -0.0999535167966372, 
    -0.113241316736061, 1.2477201366257, -0.0265419369647879, 
    -0.0935909308668847, 0.0804411654118809, -0.13974413902674, 
    -0.199298426069071, 0.118401856797298, -0.149628024097333, 
    -0.105246959487431, -0.00121575241817777, -0.0562774899459904, 
    0.035932276859492, -0.00785044556311582, -0.203185579961113, 
    0.279459534145639, 0.196899175033321, 0.234860775243126, 
    -0.122836792935186, 0.712917910331284, 0.227531641048396, 
    -0.0748437925604781, 0.241752782497266, 0.492336578467482, 
    -0.0144346070814163, -0.141854442609041, 0.12431284654033, 
    -0.0991237434722249, 0.0196328232910456, 0.000281578429866106, 
    0.0971567316837666, -0.0184701219324623, 0.106066608349591, 
    -0.179048225671407, -0.0144744256555115, 0.0166957746968462, 
    0.0288332273068576, 0.0955148321068656, 0.144206887805703, 
    0.128717356150861, 0.145166800511753, 0.0752877852228916, 
    0.0933845664162497, 0.0824739888642597, 0.0098466798563833, 
    0.0457618409830489, 0.022200097892677, 0.0286221036810262, 
    0.0254152462537242, 0.0361619342332827, 0.0431188247250132, 
    -0.00226433239260146, 0.10141825123707, 0.162160676668619, 
    -0.190924782956593, 0.0817065968989469, 0.406432470723122, 
    0.209344378539422, 0.0877319288539627, -0.0173435511918894, 
    -0.0712478974851286, 0.34552803089924, 0.113816165477549, 
    0.307307645908503, 0.783269308947287, 0.207566096749922, 
    0.0156993330343296, 0.140113170512335, -0.107325821038654, 
    0.470893924742201, 0.0297761161304765, -0.0569353105438753, 
    0.112037590866439, 0.328586324166768, -0.0188498784389591,
  -0.301030255772924, -0.0309125203352862, -0.219291661045982, 
    -0.168481679458163, -0.0760983002828863, -0.0654095434891868, 
    0.0331740667398185, -0.0953740461171608, 0.104951700966778, 
    -0.191234516814998, 0.0702050465545099, 0.0322839098287025, 
    0.0417505994919427, 0.250882978337689, 0.220916477394284, 
    0.0788548126260461, 0.0242014811047247, 0.332845518927323, 
    0.291766205385826, 0.105261672966969, -0.148176208216744, 
    0.398340294994047, 0.534584545227785, 0.146954420870826, 
    -0.282414262273361, 0.239459101191441, 0.672450931226104, 
    0.164104606809235, -0.169137946398483, 0.232521397155039, 
    0.343610765693389, 0.05731665880515, 0.649797692627343, 
    0.696783212617877, 0.405375429383183, 0.0717279450292715, 
    -0.275076781834512, -0.379115599340988, 0.683692630080105, 
    0.382058389945289, 0.0637725066633899, -0.38078885703562, 
    0.149992390848817, 0.222454505361692, 0.0238836343042584, 
    -0.0434362834762445, 0.320393104378682, 0.355016799199914, 
    -0.319861856736704, -0.236170034751862, -0.335356278845173, 
    -0.0509972889786878, -0.242520550687439, -0.0835303141323444, 
    -0.318684898123584, -0.138633721643479, -0.107834324289935, 
    -0.222969133786479, 0.156885356532781, -0.150858553225095, 
    0.224592263323669, -0.074005710949974, 0.0299275745369971, 
    -0.0578564606046959, -0.0363358985138884, 0.0232197534989395, 
    -0.061011260479531, 0.0162901896141491, -0.0301416520083629, 
    -0.0477788537722805, 0.0364761873387854, 0.0547513818907114, 
    0.0495062324234097, 0.0530597077786033, 0.0565148393531215, 
    0.0512052115590922, 0.0566328542174784, 0.0642554065085029, 
    0.0557433566424824, 0.0104156523164524, 0.286172799825153, 
    0.0834089917035236, 0.128255741067389, 0.588642509517443, 
    0.0702285935550992, -0.125855267469988, 0.081124020180165, 
    0.405339505128957, 0.142667750826735, 0.133127418717647, 
    0.214558060201312, 0.108867352930262, -0.119303035358902, 
    0.734136625293272, 0.363127606441846, 0.154256636961657, 
    0.0507150021744122, 0.345161947830896, 0.657147077606898, 
    0.0262367644275153, -0.11406510324502, -0.015040162870034, 
    -0.360396699504466, -0.0958689085847196, -0.0212715305940731, 
    -0.2543490944986, 0.0611364574951003, -0.0633868979268535, 
    0.0354436255599625, -0.255445638481709, 0.00600787207802266, 
    0.0542308057895357, 0.134592528796983, 0.251730986780018, 
    0.238958158315223, 0.17472540147209, 0.137971947171328, 
    0.176081087930257, 0.226366179405726, 0.2290444781602, 0.229715731825164, 
    0.204402891116279, 0.177065577150342, 0.201797629031689, 
    0.257861562871306, 0.247243596010389, 0.219078610746455, 
    0.253269625760028, 0.280561420783256, 0.245141866605483, 
    0.220732108239512, 0.270182514529907, 0.291811743975318, 
    0.204170918752257, 0.078355607977557, 0.199618400289658, 
    0.471551146052764, 0.233796568786884, 0.0243118838154398, 
    -0.0304088326643832, 0.550299036161246, 0.24080912789733, 
    0.0460458705523577, -0.0899986708106528, -0.0858543450737342, 
    0.414787271033768, 0.503363504641842, 0.118900900987886, 
    -0.0568363564822552, -0.176216913473573, 0.105202138570315, 
    0.641106878228095, 0.0792287089090266, -0.150805690228675, 
    0.058188672467301, 0.32310572995084, 0.084775749644835, 
    0.587742729759239, 0.316090471588514, -0.0918586235355885, 
    -0.163189536640268, -0.0701478861898772, -0.123093272695691, 
    -0.12402764922352, -0.0789122978173252, -0.159740150251806, 
    -0.067065765928627, -0.104272085504531, -0.126767748713964, 
    -0.134489542559964, -0.0235423007882146, -0.0992315854545309, 
    0.0359725811794978, -0.0298142383771635, 0.0792367052611467, 
    -0.0983880988102929, 0.0748621088695531, -0.138464324876229, 
    0.0200650272728657, -0.136067204451727, -0.0228787980969175, 
    0.0181303213653817, 0.129019747133427, 0.113991022681028, 
    0.0491308365446554, -0.0557691068168461, 0.147937336040134, 
    0.331447089692987, -0.0138138043167008, -0.253818818548209, 
    -0.265476520963431, 0.695022399360014, 0.272350544020144, 
    0.00576151839528198, -0.149107745775131, -0.0604306939753632, 
    0.855384327936425, 0.170986519733844, 0.0113821412112868, 
    -0.135257512096843, 0.456848362577229, 0.306443834290373, 
    -0.0127784017367589, 0.558448205855421, 0.259100881948145, 
    -0.305709056744162, -0.492026237126649, 0.226514044467368, 
    0.143251997081174, -0.185984238433352, -0.213458997043585, 
    0.00834906499395345, -0.231548512656869, -0.0581696424302952, 
    -0.0908628502997223, -0.0878504820438863, -0.0716812578126727, 
    0.00317951429554848, -0.181741763016543, -0.119471358735342, 
    -0.0138538367943606, 0.0547933469627432, 0.0145130082892043, 
    0.0562078814123814, -0.0166728394599676, 0.038345137473149, 
    -0.00466002836245966, 0.0332105420825161, 0.0227405913476543, 
    -0.0757106091837172, 0.144401846720087, 0.280272523902719, 
    -0.00176477539936656, -0.142041965814015, 0.423932107692247, 
    0.4715810058961, 0.121472708961124, 0.353175793556184, 0.616460020361241, 
    -0.304956736392382, 0.408827320353148, 0.754508795977182, 
    0.260740434733772, -0.440052112187954, 0.560823930535548, 
    0.882057191267821, -0.0967445563878683, -0.133622110909737, 
    0.722926697825776, -0.257691378694262, -0.348851146811001, 
    0.0171298917700842, -0.115602436180315, -0.0926408570249527, 
    -0.00121044661498892, -0.0705856727544636, 0.0608413010204779, 
    -0.159266118503401, 0.0307090862302124, -0.1301383641659, 
    0.0929649838349675, 0.103112776377585, 0.119868871916748, 
    0.252338234003706, 0.208279920605143, 0.11705601384244, 
    0.0653493890963209, 0.257212822231122, 0.208098987803987, 
    0.0838808304931291, -0.0174273031575339, 0.18908959855321, 
    0.283624709495215, 0.174655813152428, 0.151465808626034, 
    0.25804778030166, 0.270393301534926, 0.209114145034745, 
    0.193688505297036, 0.26964839767897, 0.3423139525628, 0.28777216779856, 
    0.196380165870983, 0.255642176396255, 0.387556522894236, 
    0.28820971443874, 0.141955010763733, 0.0938590481828083, 
    0.25212275007766, 0.402659522095164, 0.329877634846297, 
    0.294938880023525, 0.280683924082744, -0.136265011998466, 
    0.57820015826104, 0.236785611472577, -0.0947435778123016, 
    0.126339350023179, 0.610376198490414, 0.0799732713162345, 
    -0.0717745218660328, 0.28418964246207, 0.140092627735357, 
    -0.1937648256504, -0.119224900024869, 0.388349188123041, 
    0.180024138057385, 0.256279409057667, 0.453939616259966, 
    -0.00801723646452247, -0.110946623926159, -0.0200210882875804, 
    -0.114871323146431, -0.00544086187895509, -0.152770446307934, 
    -0.0204231558248673, -0.269908389935739, -0.0995109457154829, 
    -0.0447549621922328, -0.20621269583862, 0.0060293000367129, 
    0.0901900878141767, 0.117052154621835, 0.176425091707766, 
    0.309323394550438, 0.276776277272824, 0.122598077511256, 
    0.0325975795284784, 0.409499084182507, 0.443988828946193, 
    0.202209323387573, -0.215532285256375, 0.558258009195701, 
    0.665409569236546, 0.141149979830103, -0.396327639486455, 
    0.278184925580835, 0.596993377686274, 0.106621201594892, 
    0.0213371723945758, -0.216970644479754, 0.236311174627276, 
    0.390190809048231, 0.387123236305626, 0.250007960742522, 
    0.068002079079784, -0.172851053525454, 0.572214231244732, 
    0.255851760126419, 0.051980768886598, -0.0640016625309796, 
    -0.136693429695801, 0.0646429198905488, 0.412516697439182, 
    0.0492563798192636, -0.030196110764583, 0.00711273192415977, 
    0.368250151846538, -0.111965640836378, -0.0236119157952869,
  0.220971368928224, 0.208981992356598, 0.0553407894519159, 
    -0.0641832955692094, 0.20431181307323, 0.217261639339135, 
    0.30796384784615, 0.493067426372241, 0.25110261140372, 0.126516985761004, 
    0.154879055412953, -0.332517178101897, -0.0631606084727715, 
    0.895388576169144, 0.0528708211405689, 0.0839947123524807, 
    -0.072751633990922, 0.824306921624163, 0.00669462127492029, 
    -0.0103306432344991, -0.25532274243087, 0.345284384019609, 
    0.471264895226902, 0.0623212418262368, -0.107018831885453, 
    -0.145716091602033, 0.200478163558745, 0.387563793747536, 
    0.318612527129393, 0.162415970050258, -0.022436724802805, 
    0.331625934546312, 0.0569777026537009, -0.0497896022898716, 
    -0.0444302490677011, 0.00740476443522529, -0.145986984523504, 
    0.167597963191276, 0.219127400241707, -0.201284467984356, 
    -0.151163084191835, -0.0522471299854432, -0.110100010578855, 
    -0.100607913421203, -0.0729252297589185, -0.102359323226711, 
    -0.0252961743786095, -0.0867368596423075, 0.0550746134132585, 
    -0.138652758867136, 0.0537124003987011, 0.123563677106763, 
    0.022737671031755, 0.168788346215842, 0.194632565846224, 
    0.108856914182415, 0.347914690044448, 0.182297350600066, 
    -0.066728823026632, -0.174963476752788, 0.595891032360926, 
    0.323455275926092, 0.258589506479837, 0.1746279600485, 
    -0.425901798149087, -0.0484911021752478, 0.810724020268903, 
    0.272661610906249, -0.169120888585567, 0.320994616084537, 
    0.662273149105064, 0.305761001275569, 0.0175711188127126, 
    0.708638413187432, 0.262185119744951, 0.0507409231739214, 
    0.000886366318177081, -0.270181614729058, -0.311842633932176, 
    0.237789400207537, 0.365715559826229, 0.356921086499592, 
    0.233953242553047, 0.0915218505353757, 0.030339037507655, 
    0.135634717454548, 0.165738107688591, 0.191503091077795, 
    0.127283769002368, -0.292196775886973, 0.0668361469777742, 
    0.420129158041192, 0.139422085383105, 0.0575958251720119, 
    -0.145272217688971, 0.447324289627703, 0.294800204354038, 
    0.165362576570661, 0.0680927237264387, 0.344385562537495, 
    0.0701008829976112, -0.0896507322358489, 0.310326004358438, 
    0.705402771554601, 0.29434489075627, -0.137030418872003, 
    0.224306912975601, 0.722712432900594, 0.202240815621172, 
    0.0410736640177088, -0.0599025082308464, -0.152143949493632, 
    0.136502538093061, -0.165176963727843, 0.116053977661191, 
    -0.184257735621197, 0.0722040483011025, -0.162109552403594, 
    0.0615604189640248, -0.217657844444531, -0.0146574419391562, 
    0.105646458156757, 0.147836215299341, 0.154418388455372, 
    0.175202237764018, 0.196702644241532, 0.175464510957468, 
    0.159051408132898, 0.209339846640085, 0.211294074972502, 
    0.128405146348297, 0.0893120535314231, 0.0935410709823094, 
    0.117383455240972, 0.125223124694721, 0.101240267609927, 
    0.111590537710203, 0.129418859611604, 0.126751289725921, 
    0.105547368230992, 0.134423694951732, 0.0513492523168892, 
    0.0937882884665735, 0.359663548752789, 0.197739480327497, 
    -0.00767432512331881, 0.13157165145963, 0.390052840028506, 
    0.0846241439650116, 0.296972957739315, 0.437072894604667, 
    -0.0840398020138477, -0.0122867793251045, 0.518317294616758, 
    0.611866473968644, 0.111769531186879, -0.232003790143096, 
    -0.0573734875760233, 0.619322485755155, 0.102838176898767, 
    -0.0566694483863927, -0.0144465369915233, 0.208054139445066, 
    -0.128610829655031, 0.29599433458526, 0.287102729975368, 
    0.271362679082309, 0.362361354407025, 0.0170361438942769, 
    -0.107018025400109, 0.0198425962659231, -0.215638713353752, 
    0.142648916930502, -0.312556457656643, 0.0822472584936638, 
    -0.251022171536278, 0.0497820092992241, -0.129610912712325, 
    0.167252188401454, -0.243269692603373, 0.0954556770237596, 
    0.0413579201638635, 0.0676395606317517, 0.0311275671750192, 
    0.0762917403895309, 0.0299690816626579, 0.0529010742522093, 
    0.0782456464997022, 0.101758242899991, 0.0321117522635937, 
    0.0811057218590055, 0.103577733863606, 0.10865038494446, 
    0.128944064300809, 0.138235992699801, 0.121388445437683, 
    0.139976096417802, 0.12778749597396, 0.000725335498636209, 
    0.158766184188563, 0.32532873367853, 0.0572526168215815, 
    0.332823502632454, 0.455723773271753, 0.125821751592265, 
    0.0108009053956906, 0.537714083596387, 0.321365200578762, 
    0.0953572230473035, 0.195520146727045, 0.493991541723071, 
    -0.092558710041519, -0.311108217671701, -0.303011008818567, 
    0.470607346547787, 0.439491780623369, 0.326152552459405, 
    0.521285547117008, 0.158099291343149, -0.42208682596052, 
    -0.233940105577468, -0.203674153519858, 0.00608285004112297, 
    -0.214492386607148, 0.308676392943042, -0.28381163961249, 
    0.0224835846819978, -0.190753325208159, -0.056101112663915, 
    -0.315890315239362, -0.0499195905997977, 0.027275132706382, 
    0.198823988393529, 0.252236569152846, 0.228817578628102, 
    0.185511876292474, 0.201417191038768, 0.321501708052771, 
    0.35187632545004, 0.24250514544025, 0.151310494025799, 0.140157697598501, 
    0.113392015995729, 0.136059905258044, 0.109137472061931, 
    0.117467307818393, 0.105304197194432, 0.145268905922528, 
    0.146231046243075, 0.0554072034078333, 0.543472990931384, 
    0.0556911391337787, -0.127834396994785, -0.148903223379146, 
    0.539854849301853, 0.324553034572127, 0.0920869197224922, 
    -0.0924027105693706, -0.0161036950433344, 0.354807114920156, 
    0.303091444555148, 0.18191275376865, 0.0574001761825777, 
    0.186445269008167, 0.337418216900337, 0.131243970890988, 
    0.0528258458206868, 0.300385260250917, 0.101424849074145, 
    -0.0364918576268977, -0.05349948240218, -0.168316870322858, 
    0.0841657326455584, -0.132957866588275, 0.0502610110736956, 
    -0.161877994972073, 0.0356178034750748, -0.112622117705659, 
    0.0557393360024718, -0.233111605731391, 0.00853440176371965, 
    -0.0742291870617679, -0.0557186673162419, -0.0614028004416164, 
    -0.0520204723921036, -0.0594046777373512, -0.0319758312653434, 
    -0.052469696222442, 0.0521732519394728, 0.0318278664239166, 
    0.408823061431407, -0.34664401486061, 0.0451434856282442, 
    0.770019860504481, 0.613089872743631, 0.264690398374799, 
    -0.0202809810970061, -0.162559359025034, -0.269506308946744, 
    0.418692542661406, 0.314227116299341, 0.139981562225305, 
    0.344273733566692, 0.494530165790892, 0.223343878041607, 
    -0.392122715663013, 0.373458453777013, 0.542402950946141, 
    0.157763302410928, 0.146043049818037, 0.495330903978718, 
    0.0341430321377433, -0.0779536685042334, -0.10377761413054, 
    -0.00711313069947511, 0.0571201661564859, -0.0498903995454018, 
    -0.0479675917938535, -0.0302204093732211, -0.0667654536048695, 
    -0.0156638304811001, 0.0606327837911837, 0.261108749146203, 
    0.194691195240958, 0.0571628655436861, 0.34150434043652, 
    0.43004350705701, 0.144352165399512, 0.078722448805941, 
    0.155448993930934, -0.245308146580027, -0.108537520063003, 
    0.796914259422296, 0.433436047948253, 0.165289136888068, 
    -0.182357380862111, 0.282487210467756, -0.144940763427853, 
    0.530848873725447, 1.01163373102146, -0.0288973075145278, 
    -0.119970002720865, 0.316984995297208, -0.271212979217686, 
    0.507476816094045, 0.130951353841612, -0.0204403390581184, 
    0.346431291328478, 0.0658672657030281, -0.130849581312944, 
    -0.202504730122551, -0.0944740638817865, -0.223283029794813, 
    -0.138734431805844, -0.113774483962321, -0.179080325526361, 
    0.00663046292502481, -0.079524742370503, 0.216816836376261, 
    -0.195360573815141,
  -0.263148397953979, -0.124469573324055, -0.340656706386789, 
    -0.250922781144193, 0.157585308665903, -0.230575441038937, 
    0.100016047474446, -0.0642649549204031, 0.0680461878721968, 
    -0.254031896668873, 0.0063681455747204, 0.118606103764703, 
    0.138889223420879, 0.145683357786249, 0.1426305003077, 0.120960894884173, 
    0.152285070497772, 0.205569679837353, 0.15955458635912, 
    0.0911830932076994, 0.128418664705414, 0.172792259497468, 
    0.149340867920187, 0.102833541606001, 0.223156132377911, 
    0.25727974670294, 0.120908703537705, -0.0166935398645783, 
    0.129730793650233, 0.265436507575239, 0.0717421141028115, 
    0.361541411078692, 0.823553195637754, 0.235316901193365, 
    0.235792565931934, -0.108319131800016, 0.723985758818225, 
    0.0926194049221298, -0.153225009811527, 0.0239166199786081, 
    0.448416161047409, 0.211781338507632, 0.00282151994488955, 
    -0.111479653435351, 0.0271057036273316, -0.060785126305515, 
    0.306363669503915, 0.142443530403729, -0.0156910037185083, 
    0.00676338274148509, 0.0139284659835506, -0.0977689282498583, 
    0.218468486074967, -0.045503861567638, 0.21782559660329, 
    -0.188557842036732, 0.14497308610966, -0.164168565374063, 
    0.0995283996424909, -0.292207923468756, -0.0238730240191551, 
    0.0694595922271691, 0.112577982549669, 0.163905237977456, 
    0.233167793857168, 0.221237809890956, 0.146942802231284, 
    0.145704961941114, 0.280455562518483, 0.259608837880069, 
    0.162758789975979, 0.135738389757307, 0.123817143240478, 
    0.131729783794045, 0.138946745536042, 0.111771372464979, 
    0.102629190897114, 0.145240017513249, 0.154956696656723, 
    0.112104594688811, 0.103217284869812, 0.102798931801394, 
    0.124643197645007, 0.225133348709976, 0.217603952650912, 
    0.118891313879486, 0.081834486495878, 0.19926639271572, 0.14291436965203, 
    0.0564975682531504, 0.435050792161841, 0.404725111778428, 
    0.196210612176704, -0.135489455957785, 0.667058686993189, 
    0.342572328789439, -0.250928278035839, 0.686016569227333, 
    0.540419959456303, 0.0776108372487749, -0.158328286880925, 
    0.219487963120191, -0.114217829174036, 0.173103852069665, 
    -0.316018099622197, 0.0285289299750982, -0.320209176415678, 
    -0.213527288277941, 0.0867666111097324, -0.193370767815902, 
    0.216151207477083, -0.0477251756856088, 0.018297021777518, 
    0.0761745152545224, 0.0733756841444788, -0.0720826091440549, 
    0.0403410952572885, 0.061448977761279, 0.0904118804666763, 
    0.00769482665056065, 0.00501758823393856, -0.108877240162466, 
    -0.0262991612436992, -0.0688687854853772, -0.0360131869387761, 
    -0.0622617011213253, -0.0209714091227012, 0.00981835679577681, 
    0.0777783166483866, -0.124857575479421, -0.0680848116059807, 
    0.155179535526137, 0.251294957492055, 0.163070087632889, 
    0.0805676806509715, -0.19194361660464, 0.151456190862475, 
    0.349268754733122, 0.116557268882821, -0.000486214214971886, 
    0.191297851654724, -0.00600101191696653, 0.94869267665708, 
    0.462845026567075, 0.0811407485187575, 0.315598364602747, 
    0.634251528641412, -0.0490188783422364, 0.552114312837051, 
    0.873530558108264, 0.0838481185796509, 0.061149049563698, 
    -0.155729414123294, -0.00943439254684375, 0.184499746947085, 
    0.478967764744721, 0.201048266705312, -0.115966570607165, 
    0.284007770551496, 0.218986651658476, -0.199416515579358, 
    -0.0378329845240572, -0.169057407211284, -0.0826097959630124, 
    -0.021920999904607, -0.174958939528018, -0.0943874608433147, 
    -0.0684870568387982, -0.0233534303071919, -0.0883527358793772, 
    -0.0346359717248741, 0.0423943446664644, -0.0786677320661836, 
    -0.00756315237035518, -0.00806862269169681, -0.0438124837687266, 
    0.0211716626748385, 0.00551868538479198, 0.0384077337843894, 
    -0.0543960806172133, -0.0233554011495751, 0.199503887062272, 
    0.167804049078353, 0.0310112370026097, 0.00245861194898146, 
    0.27685051709508, 0.308047790328613, 0.216997825472878, 
    0.154480700583685, -0.341853221222648, 0.173067886426352, 
    0.41220161043663, 0.318849539876045, 0.498913467422075, 0.28743363326916, 
    -0.297011392670761, 0.0551863185065074, 0.586662445338843, 
    0.369388286965828, 0.126679859780175, -0.201650818563102, 
    -0.0522229542385237, 0.314774535742848, 0.402745596532697, 
    0.0876554296295804, -0.0723168604551195, -0.0917711473865052, 
    0.330130659976078, 0.0331553034029432, -0.0553639271276141, 
    -0.314699445818003, -0.0390099973530948, -0.173357080989415, 
    -0.239507408602194, 0.146089817819395, -0.201498431844778, 
    0.039054982097421, -0.124877698351682, 0.0131413812935101, 
    -0.259231648556032, -0.0314378882147647, 0.0582317358783251, 
    0.0997615678353514, 0.160409387095712, 0.184788060145297, 
    0.143078949517156, 0.168319982053238, 0.23469612418001, 
    0.141676399262552, 0.0984498807094204, 0.412757612976318, 
    0.262057228599418, -0.0332444894493186, 0.506401550827082, 
    0.54030889873362, 0.192478043797067, 0.0786767186673949, 
    -0.124648330793377, 0.249629962399087, 0.741711836163002, 
    0.357031838586507, -0.00242288952663682, -0.240597926154993, 
    -0.16914100213775, 0.497615917840496, 0.240994297188142, 
    0.174415847177711, 0.221373235949856, -0.189999576490191, 
    0.406470555247824, 0.265370510744043, -0.102340367891403, 
    -0.12570611900565, 0.0213347441236006, -0.00453028649025308, 
    0.168067964595606, -0.0886428005507717, -0.115500096675557, 
    0.0223613801475523, 0.110625341890498, -0.0252630906256858, 
    0.0140138901060677, -0.0457892663875554, 0.01634913713661, 
    -0.0706703535189747, -0.00642608127200434, -0.0305418748659653, 
    -0.0177181443869092, 0.0373029056945646, 0.0226789598445605, 
    -0.066739132164122, 0.125911525882297, 0.216042883978642, 
    -0.0611669689256598, 0.358579456153999, 0.569050716986157, 
    0.11556985014321, -0.186574429641877, 0.0330117202952744, 
    0.461441872416604, 0.369280730100657, 0.22235704688488, 
    0.408931834844017, 0.168416372447896, 1.21315638319141, 
    0.380136520642399, 0.0371841070467301, 0.488201160275214, 
    -0.066944377987609, 0.689640020656313, 0.13234916908752, 
    -0.02167595990869, -0.104045952881262, 0.0330950677690719, 
    -0.00305884125697048, -0.0412118611104339, -0.0442927392132897, 
    -0.00934275788285957, 0.0706226257373725, -0.10111420723184, 
    -0.00730253206378742, 0.0148072924181156, 0.063380859597289, 
    0.0299981268955992, 0.0398993466432115, 0.057458753618176, 
    0.0978121465564974, 0.00599918722958967, 0.004358611085862, 
    0.0605599952302106, 0.0295597179387264, 0.0496971812248488, 
    -0.0362171023252212, 0.0258217720501239, -0.0635081695394327, 
    -0.0337009074409244, 0.0301225015243983, -0.0147666993660282, 
    0.0612197980298511, -0.0274183689886723, 0.0531299148078153, 
    0.0397565329010832, 0.0513427594198318, 0.0520691274760318, 
    0.0606484190513365, 0.0264272403391578, 0.0443746085918283, 
    0.053898756246222, 0.064067233039972, -0.00653903121586257, 
    0.0999856363495592, 0.136528532084198, 0.0761130757142584, 
    0.128714198011811, 0.267937678556054, 0.180032302863196, 
    0.076396347214637, 0.133178920064409, 0.169569398499848, 
    0.136567747953811, 0.395820378378138, 0.375884755500474, 
    0.0725344711863742, -0.14880463962823, -0.163691024156369, 
    0.360142891970742, 0.462849067392041, 0.198035833551028, 
    0.242949534895845, 0.631248526684685, 0.292202773388275, 
    0.190713265169198, 0.0512851671768301, -0.163529891930501, 
    -0.045001803875096, 0.122809546808012, -0.0674105813668715, 
    0.301866534073361, 0.275665527211121, -0.113268854470035,
  -0.0550816204050159, -0.166667207144861, 0.21557475243787, 
    0.29446053181844, 0.44007574219779, 0.0172972135279942, 
    -0.123871226777857, -0.152337091542171, 0.0794711959021987, 
    0.253247102914774, -0.119217248133687, -0.0438720846128662, 
    0.00165082755654138, -0.0513889550663137, -0.0483832440901298, 
    -0.0278701214828045, -0.049697592984363, -0.0193862574808033, 
    -0.0208825127352094, -0.0975196372641523, 0.170661373623778, 
    0.113810407518618, 0.0147784530459859, 0.256934643757353, 
    0.176036317563792, -0.0324399960614104, 0.394945476851956, 
    0.452493820119557, 0.0304579474795659, -0.197766887829588, 
    -0.00432949367986746, -0.0172115409468922, 1.0022796202259, 
    0.279440164694857, -0.0878508550253912, -0.028949702499664, 
    0.018428806877842, -0.216265148457232, 0.978398181633436, 
    0.204100098427257, -0.0905245959977326, -0.210528058581628, 
    -0.00339188434338794, 0.0785163172130731, -0.100446006095762, 
    -0.0273275686073803, -0.077092312104125, 0.106084155074353, 
    -0.0161135468876951, -0.00746281862038365, 0.00324486539844243, 
    0.0665437033672369, 0.0290858511649447, 0.0212327312610333, 
    0.0336613069593797, 0.0491794542165553, -0.079525471176879, 
    0.13758642031058, 0.232613595170074, -0.139580267447452, 
    0.128538443330917, 0.26098658620441, 0.152728222403916, 
    0.593712519256295, 0.491607228279579, 0.206818866222624, 
    0.495695411979295, 0.416391927239298, -0.338708044263293, 
    0.307960398935498, 0.713590882279422, 0.524938930081978, 
    0.59979609751736, 0.34003551262538, -0.193626216570869, 
    0.413471534859527, 0.340437642763363, 0.44640491822698, 
    0.602631727954999, -0.236485691021457, -0.388888826291032, 
    -0.038701057581715, -0.134680111281247, -0.163035928592035, 
    -0.0789879076558998, -0.161145870760256, -0.0548927879666343, 
    -0.113254001015048, 0.0495095365320004, -0.221461437763926, 
    -0.0931919076400738, 0.260518914993421, 0.257120375438404, 
    0.130931360171158, -0.136027792307572, 0.361958753922476, 
    0.403012726114398, 0.140145825145049, -0.0810784146194843, 
    0.293445465882649, 0.338531944287877, 0.184139112979698, 
    0.118459374043028, 0.114481088210203, 0.122719579705222, 
    0.130294525598494, 0.124411048890954, 0.12434478193443, 
    0.0757344374070526, 0.0672564499511407, 0.0894259133680492, 
    0.114549425793028, 0.112968819320046, 0.115271364105959, 
    0.167144402301095, 0.2016427357786, 0.170530179056057, 0.111016837730229, 
    0.078099797586678, 0.321808467379154, 0.276357661659277, 
    -0.0363058821079336, 0.0195358945647143, 0.501546546937096, 
    0.334727305633895, 0.215762332509293, 0.149091958663804, 
    -0.104233737609143, -0.0302952836617774, 0.75433240545863, 
    0.148239397902074, -0.0628397040838133, -0.07723465265858, 
    0.0759523985536716, 0.331557350392633, 1.03457449231705, 
    0.368536082238436, -0.0411354531459535, 0.385385885681552, 
    0.485193630828825, -0.124139679125859, 0.113102825334966, 
    -0.416814782938197, -0.0173798809963786, -0.350335042511124, 
    -0.234777381595048, 0.00803508960176512, -0.258269929914022, 
    0.135009690801682, -0.199742762104658, 0.151527430144994, 
    0.024555692236023, 0.070148227580258, 0.00918267732524881, 
    0.0528540313016328, 0.0308171323625644, 0.0657461216264658, 
    0.0573833939089896, 0.0529675407030084, -0.0830758915239485, 
    0.0143666332035225, 0.0882260404976975, 0.154212778600522, 
    0.126492556407149, 0.0623079679597867, 0.134376152774112, 
    0.282336992253257, 0.240895410748889, 0.128408895009698, 
    0.0493296307957959, 0.169970076529074, 0.291699268540019, 
    0.247558691183582, 0.217281786806077, 0.331164044732438, 
    0.37842521787797, 0.255608222341961, 0.12170540589762, 0.112858239353453, 
    0.418293505931663, 0.420779895068844, 0.155459976432737, 
    -0.121155465596494, 0.275636821861574, 0.46761234431294, 
    0.167117982844831, 0.0885286858740295, 0.630422185370268, 
    0.219569243178962, 0.0135460686446565, 0.571464103808198, 
    0.105872477559244, -0.0587277715441376, -0.320423761697982, 
    0.152951814154696, 0.600598118434214, 0.28280421386818, 
    -0.124440160913086, 0.25824874671988, 0.406132168377534, 
    0.113313550996377, 0.0269916703334659, -0.18397853584561, 
    -0.0676591613711259, 0.141663104505227, 0.0814105941798324, 
    0.0768708225615841, 0.0850196419608729, -0.115162702843998, 
    -0.234890540410791, -0.227878335240018, -0.069432373191453, 
    -0.256094808915032, -0.0875684200077547, -0.227912483295029, 
    -0.1130457723947, -0.174284896949654, -0.165272578832958, 
    0.0397302424547782, -0.204426451587417, 0.115194820796035, 
    -0.0515215625057671, 0.0217167138264602, -0.0349249869286081, 
    -0.000389094895687878, -0.00346082413168317, 0.032902461513154, 
    0.0171297169735257, 0.0652885875374551, -0.0760255095968177, 
    0.0613382627944667, 0.0609717923940155, 0.0156373886901384, 
    0.126224227457274, 0.17056975172366, 0.0839599898815998, 
    -0.0452137471925235, 0.152719809773417, 0.271668408337475, 
    -0.0670604428439599, -0.127650069076941, -0.391497563565841, 
    0.654984646995449, 0.294091376181453, 0.101957403532241, 
    -0.304427084574146, 0.321452104732725, 0.487271888520094, 
    0.289106373206662, 0.444972868986298, 0.358474731505928, 
    -0.00376358064024868, -0.0139039290096894, 0.0137451611591862, 
    0.112629801135439, 0.250017891739986, -0.0513737786040452, 
    -0.0215039628428956, -0.0381421509571565, -0.208267688401434, 
    -0.329419377816843, -0.0503159313106683, -0.268437067630062, 
    -0.188636381114016, -0.0994183724300408, -0.191876793127769, 
    0.0331450303565702, -0.210306416598307, 0.0661698840298139, 
    -0.1244435904839, 0.118586462445794, -0.0259963384049087, 
    0.0305023956471751, 0.00844818669736776, 0.0400995069960869, 
    -0.000535261613916205, 0.0504670923862284, -0.00856311093047023, 
    0.0441715193800146, -0.0469443963943613, 0.0557026207769232, 
    0.0406815782867495, 0.0518246805417022, 0.19815568606412, 
    0.124454050743679, 0.0320704171459163, 0.0370769706646222, 
    0.13468058679844, 0.0905254075587176, -0.0309319714285864, 
    0.489498513484712, 0.358387335814651, -0.0127542930077512, 
    0.0808236084366097, 0.700614470238507, 0.878670544618011, 
    0.0134660465511023, -0.308113133079919, -0.182337049110918, 
    0.530353231893034, 0.193005692470617, 0.0504646511892363, 
    -0.184893396322968, 0.0581718885873701, 0.142747289933624, 
    -0.00764571293300653, -0.111691295332958, 0.198609714421592, 
    0.131892032585243, 0.0366203595931727, -0.122860154590168, 
    0.109898523076448, -0.0812504880683481, 0.0649133711295902, 
    -0.403456606827463, -0.0200092282827306, -0.118478955650501, 
    -0.0892093965609675, 0.0497857129987729, -0.306374584183205, 
    -0.0565298990307085, 0.152158790069329, 0.0226438497817431, 
    -0.165692625969343, 0.189621354209178, 0.315556830070674, 
    0.0205527619659406, -0.121103140456262, -0.0914789268708306, 
    0.203405740623098, 0.147874939239702, 0.668996429543257, 
    0.792412143050668, -0.502594504545024, -0.430283800168154, 
    -0.253987325883132, 0.807426019237991, 0.235213915777701, 
    0.264558593689109, -0.057673548566603, 0.723215240038431, 
    0.339378913609159, 0.194641985080864, -0.25725899205234, 
    0.335786963130672, 0.533934948576158, 0.0765523403262375, 
    -0.193172076538062, -0.0563249493684146, 0.569787124686713, 
    0.124190813348901, 0.134564958033105, 0.331983612912585, 
    -0.0535483572220211, 0.547130140630106, 0.226766846053639, 
    -0.105797860257049, 0.284711748319838, 0.328338969466285, 
    -0.13066692904357,
  0.0396016012612192, 0.0819095401633609, -0.151674999730239, 
    0.221916380553984, 0.186082605886526, 0.0420363375161937, 
    0.494387085506102, 0.178260527872072, -0.181823794709169, 
    -0.0717028169243433, -0.321113276686796, -0.228132964167322, 
    0.0568379926052795, -0.187522524489915, 0.147497566334742, 
    -0.280372883676477, -0.00139573623885562, -0.0875395814270149, 
    0.0501550985793478, -0.287623446835143, -0.00360309739498488, 
    0.0828001499944805, 0.0974931404778048, 0.149699997301995, 
    0.177183949914212, 0.122499182238423, 0.110329268630513, 
    0.177081715127486, 0.159215567835566, 0.100675702748352, 
    0.142056108348094, 0.146867827498588, 0.152869365568818, 
    0.238380568050236, 0.247449856217768, 0.129174987492956, 
    0.186764620968239, 0.443859394576382, 0.184352037466137, 
    -0.0597020920016996, 0.0357485026173755, 0.574948698453974, 
    0.14880669271635, -0.046250075174331, 0.0032793530405418, 
    0.141421472729401, 0.367819145132787, 0.64028532116467, 
    0.262306794816554, 0.0419756320444687, -0.402538917177683, 
    0.308860834366344, 0.485342901712747, 0.117574709445511, 
    0.015915781706319, -0.220743170675712, 0.0366227944669743, 
    0.161937208615267, 0.684211829068491, 0.281097916872449, 
    -0.228094331824441, -0.152548212302868, -0.0917886498719218, 
    -0.129270049005916, 0.112787761340238, -0.120037253405882, 
    0.0429382841763272, 0.0496146617544657, -0.0197927489650704, 
    0.0553463996308455, -0.365575271299967, 0.080060947821801, 
    -0.181148259901078, -0.169131577541653, 0.123348871069875, 
    -0.16162349090959, 0.0541135109972575, -0.110096350411585, 
    0.0533087263447562, -0.385843477105567, -0.0206728905047521, 
    -0.0244332730499132, 0.0223496705444528, 0.109555430456878, 
    0.0447031527374121, -0.137038142073343, 0.114025937190689, 
    0.161036239779916, -0.118922345332235, 0.00170522755208263, 
    -0.0422175307064591, -0.158637956243773, -0.0933924751376707, 
    0.419374610576322, 0.777388973790792, 0.166181853359004, 
    -0.270093915864957, 0.173482048091723, 0.514850120832932, 
    -0.0979409844055139, 0.322347697161462, 0.935234704336981, 
    -0.0720359498977648, -0.0937375690354188, -0.253391598782423, 
    0.82854610911739, 0.231061866023776, 0.0041117002299659, 
    -0.0746125270852778, 0.381636581562057, 0.515041055143106, 
    0.29037070597601, 0.00740030296115681, -0.104053931710947, 
    0.843174960195013, 0.296400026198977, -0.0032305547241441, 
    -0.313271264555911, 0.0855101483944355, 0.533652640553108, 
    -0.0947527966471808, -0.13726516782358, -0.00995277057167802, 
    0.305316044787463, 0.0564353605127506, -0.151271460972467, 
    0.241909957786855, 0.318235863987144, -0.00822720462876289, 
    0.282122529911267, 0.0272605154739762, -0.230671806200186, 
    -0.165034645034487, -0.0972900911320943, -0.161271464354564, 
    0.0423864080446084, -0.138912663900631, -0.138277140921463, 
    -0.00599603629471382, -0.0610691743776715, -0.0498664151593705, 
    0.079942017844071, -0.137416520842596, 0.0220310201928573, 
    -0.11096347148917, -0.0318726895686467, -0.0717787952548785, 
    0.00104012099674955, -0.0846212488609705, 0.0192923945632704, 
    0.207928349307534, -0.0574841290753499, 0.312923532426696, 
    0.260556742138317, 0.0499236646273715, -0.0121960259578489, 
    0.435643015823502, 0.177069731860326, 0.0246613397193003, 
    0.015417169660539, 0.301047470486832, 0.0387741365435661, 
    0.501105824513258, 0.584092291795878, 0.276810316405246, 
    0.252455305446603, -0.0532887951205255, 0.724210499555857, 
    0.606262736255225, -0.0614590586965078, -0.172372105687135, 
    -0.000646015218736001, -0.178757498605274, -0.0951635645500403, 
    -0.00287919971027938, -0.164471308955026, 0.00852592894675358, 
    -0.0490930914436288, 0.00376517444629798, -0.136108654741491, 
    -0.0136134405329733, 0.123612037906537, 0.162012780601993, 
    0.119706774681323, 0.163881354541469, 0.301349332297937, 0.3122774716971, 
    0.169083587019154, -0.0152577345842121, 0.371543875637361, 
    0.619487525193867, 0.265529712783546, -0.241377165030566, 
    0.720819269896589, 0.432215398932103, -0.024371416143892, 
    0.518256081199472, 0.587928634896192, 0.15405801866783, 
    0.0401995418401387, 0.592416418148767, 0.993940431416883, 
    0.40234874382442, -0.178820832601892, 0.612793222605921, 
    0.538602332760287, -0.000626910154610957, 0.660317218763206, 
    0.728658743897049, 0.0681530549567122, -0.0161510230568948, 
    -0.13416525726893, 0.0819342709958496, -0.0944879704353594, 
    0.0650619059954109, -0.201650617564396, 0.509686963518267, 
    0.491942551314167, 0.113169868371396, 0.0525405877188771, 
    -0.136746372041327, 0.127918743193939, 0.0327516579456117, 
    0.0872586716294813, 0.005073245275853, -0.0102433866770835, 
    0.00102768456444852, 0.0361838172959448, 0.0384747435991422, 
    -0.0340796507631518, 0.51230747901249, -0.00688548704586775, 
    -0.0410572147523084, -0.271313972606597, 0.460460235228692, 
    0.399192739184587, 0.0779969266269736, 0.448463119705507, 
    0.525516940257956, -0.0328672741157927, 0.340543821924169, 
    0.618873942127309, -0.470381748349265, 0.229104594796114, 
    0.693589358247283, -0.11714784680218, -0.474956289119645, 
    0.441065123819447, 0.492939826071435, -0.416771684613435, 
    -0.0936830933225134, -0.136916324958964, -0.0627448153387698, 
    0.270132191022557, 0.101581712465548, -0.0854124485232061, 
    0.111515366153503, 0.095524275909888, -0.034582906626856, 
    0.0337983200112546, 0.187278307993794, 0.051390693107225, 
    0.0203939379664468, -0.0589203678219438, 0.0581177222734315, 
    0.0953838169931365, -0.0722795276957262, -0.0853463043445866, 
    0.0715741994831271, -0.020336320199142, -0.136685887304354, 
    0.0527080017421274, -0.137662864922041, -0.0403793867410222, 
    -0.0430442143165486, -0.068955604538119, 0.0644573299020339, 
    -0.0783641994194938, 0.0872459743774603, -0.0696160667091121, 
    0.0608827849024366, -0.0679197046955998, 0.0159094738890036, 
    -0.0298341018446546, -0.00453211318895741, -0.0912371110788672, 
    -0.0300687624112375, -0.0204248854523165, -0.0846659083618193, 
    0.0148814144616345, 0.00820502028374719, 0.0829318340692442, 
    0.12460762734338, 0.0847298378130945, 0.0572172092512639, 
    -0.0642303279762016, 0.0918657807519927, 0.276233020815329, 
    0.0413902732169698, 0.000110763096114519, 0.437838338239448, 
    0.443854089739392, 0.5631360921365, -0.251034532820559, 
    0.755365491364423, 0.524939543906549, 0.121428832598138, 
    0.180872705893668, 1.02276146925383, 0.302299007457406, 
    0.0308267863187713, 0.0393213045464871, 0.0584805935526269, 
    0.0984161776596018, 0.100612907604349, 0.0921479665186725, 
    0.111289461297163, 0.12093708779434, 0.103534395916126, 
    0.0737198967416243, 0.0670977319055506, 0.0740434772235937, 
    0.106567615063, 0.150272181574207, 0.134437068265595, 0.0877491882780683, 
    0.0875227267917843, 0.160014294839122, 0.14166710764196, 
    0.0727242010779512, 0.0615726447025768, 0.097109871385116, 
    0.335016877085477, 0.316203428482887, 0.121202949802881, 
    -0.0402769508346092, 0.00407852357321521, 0.414375043858019, 
    0.364778704138147, 0.165617353121352, 0.0662494231571593, 
    -0.0613583306643071, 0.440444902914637, 0.409620871914437, 
    0.120899865908701, -0.0623885817323264, 0.542316024993728, 
    0.399600910885624, 0.116862303799765, -0.0677125713809694, 
    0.573596049061725, 0.387410616914562, 0.104631465560747, 
    -0.228684427948057, -0.0306708612488156, 0.559572047425485, 
    0.112888961737318, -0.0619578877240079, 0.0827439868489281, 
    0.514143445861894,
  -0.326326417852264, 0.0186708977739933, -0.139227269949615, 
    -0.0346111109044648, -0.194321998032348, -0.121329238249608, 
    -0.145725223832468, -0.123587627800656, -0.116774479681052, 
    -0.12334168977429, 0.0570268611972717, 0.0702364928495033, 
    0.065974759034719, 0.0851324082451904, 0.078962425064533, 
    0.0485255889534258, 0.0425244103329085, 0.0515370781452194, 
    0.0484118644553726, 0.0540307110351077, 0.057797182650087, 
    0.0108970515123557, 0.0485430752527134, 0.0578243443172032, 
    0.0590366234526058, 0.0281292902802318, 0.0442495998288122, 
    0.0609868153166616, 0.0721300001608885, -0.0108432131501772, 
    0.119586892216774, 0.152120889230475, 0.0617391999820739, 
    0.151610662159499, 0.243791455160014, 0.0923540887002692, 
    0.247869297644568, 0.370150235707814, 0.0692569700857459, 
    0.0606256399499288, 0.196275517495517, -0.291656990092954, 
    0.569162373557507, 0.328812040020981, -0.0318283361033529, 
    0.310731523318849, 0.430243463888158, 0.0934462087419443, 
    0.707054909031312, 0.357755308169889, -0.207313115598585, 
    -0.129792467655364, -0.15486880405932, 0.0783917694819012, 
    0.429126594737042, 0.160225980361584, -0.106699464986511, 
    0.181076633408718, 0.374783042807565, -0.0497171591880988, 
    -0.0533856742604593, -0.145704746480649, 0.0775712815466556, 
    -0.217765251340129, -0.0355068325155715, -0.253258564343719, 
    -0.145097630695029, -0.0904462760155483, -0.156175570288511, 
    -0.124198109590575, -0.133234653143321, -0.0427830509549241, 
    0.310096841170582, 0.239443182629819, 0.0377806734559395, 
    -0.0782148917726471, -0.205991561563154, 0.449507105426396, 
    0.270203352381921, 0.203739313858183, 0.0382233497578818, 
    0.91070707666864, -0.0938175754000282, -0.52187065669467, 
    0.159564443839022, 0.620207565588702, -0.101730198546074, 
    -0.0825746762108242, 0.0724454968427444, 0.810264707859585, 
    -0.0929341951674193, -0.000484299552379067, -0.0318579526203668, 
    -0.138399632201787, 0.427077650842585, 0.344696485090331, 
    -0.0535700307409191, 0.591055533291832, 0.374213953047357, 
    -0.119566480282174, -0.133605649294558, 0.0743403087280573, 
    0.00315817897699842, 0.211271323931926, -0.0751585671361087, 
    -0.00849803671864699, -0.0841832342123234, 0.118437106142376, 
    0.0403734357292897, -0.0173554070943133, 0.00208074895241192, 
    0.0735460272904896, 0.176810696430127, 0.19991277208219, 
    0.142697655199664, 0.0897529632447145, 0.092079987860827, 
    0.121938931906019, 0.190496618308973, 0.16162871293227, 
    -0.125121200471056, 0.295844651497837, 0.466980958148681, 
    0.168493629630759, 0.0379260921034887, -0.0315554844826371, 
    -0.193900841466825, 0.313672054201786, 0.429688933154757, 
    0.320581604495411, 0.227888783562654, 0.104690246883135, 
    -0.0922444843423187, 0.476833817796456, 0.259967417124635, 
    0.0621086092384707, -0.0213687411895398, 0.390520466538591, 
    0.169379710745495, -0.00917216425939089, -0.0872089890278546, 
    -0.186591366207955, 0.047722966233047, -0.079864773843737, 
    0.0365567132994423, -0.155338268833563, 0.0368178212665174, 
    -0.127160020798983, 0.0157029701044263, -0.174054295669177, 
    0.0038985430279599, 0.0911938056551856, 0.014279083552936, 
    0.196455552550461, 0.392707002496472, 0.0753429530369437, 
    -0.157506148485375, 0.023854725402129, 0.437913304924579, 
    0.155402954838998, 0.230676058322345, -0.280739037354315, 
    0.203669065651395, 0.65653660541541, 0.213078786454683, 
    -0.153912433139966, -0.0417508049573753, 0.46787584818011, 
    0.57217327357344, 0.200839861031306, -0.206902299058049, 
    0.141241353942193, 0.359521856957503, 0.105792010686848, 
    0.0649435649729873, -0.174139964583807, -0.0199757378579669, 
    0.152002789860476, 0.31799796833342, 0.220354198048924, 
    -0.0893696373669702, -0.129726604792498, -0.143032014119445, 
    -0.0815673624710839, -0.00149024899240881, -0.1830536050804, 
    -0.0805310402201705, -0.141770268944246, -0.100865962211439, 
    0.0272673068416654, -0.119987101683747, 0.103482628577313, 
    -0.197060237066517, -0.0629643383512516, -0.00396478375415346, 
    0.0558103040489072, -0.206114812832108, 0.0543204178353714, 
    -0.293619447748544, -0.162940447443717, -0.0353340360382409, 
    0.0745564362074242, 0.0551505985697008, -0.000415777395235434, 
    0.188412915912289, 0.151023501071858, 0.0209393842398143, 
    0.0406586958017474, 0.130124146889885, 0.362317372428055, 
    0.271962027091877, -0.133771881652145, -0.103809833224263, 
    0.73996614608779, 0.151384669166453, -0.0586603002420938, 
    -0.197852349123029, 0.173128938420823, 0.746105507403979, 
    0.318437910491342, -0.109801665501885, 0.35087076203507, 
    0.412398073576914, 0.324777680302629, 0.245796088463313, 
    -0.32885959632809, 0.172412228121948, 0.330928624208336, 
    0.470211557171806, 0.701651799472891, 0.0910471492843781, 
    -0.111189998868263, -0.168314890509325, 0.19532382232007, 
    -0.127522355300795, -0.0525617309864072, -0.151810398253858, 
    0.0483973029387768, 0.132415980357336, -0.138316969065191, 
    -0.029941522611774, -0.055669244988099, -0.0363309937536356, 
    -0.0523510815424205, -0.0469860537706604, -0.0450444173341528, 
    -0.0460322974339285, -0.0321078576867872, -0.0438235469319224, 
    -0.00342916722589816, 0.0925728604381087, -0.056602479488408, 
    0.152200899805434, 0.309329531649859, 0.156294535680133, 
    -0.0602283244414505, 0.268520020859614, 0.438968424774549, 
    -0.0622574211929695, -0.376600142446155, -0.154020015638404, 
    0.634321604254224, 0.0942797619494037, -0.0190996300033514, 
    0.325879216306015, 0.262575752629414, 0.0827176650549784, 
    -0.54585047148777, 0.453746664007541, 0.0101036782685004, 
    -0.38478119498591, 0.0921934964021235, -0.125880268326393, 
    0.0775485371897062, 0.0539665482156178, 0.127762046510484, 
    -0.116829714384625, -0.138006166555777, -0.229236791114639, 
    0.0387100552420117, -0.292910608618134, -0.0686892665634447, 
    -0.0590303012510115, -0.174537434129428, 0.151157224277925, 
    -0.214011411661907, -0.0061342272667944, -0.0160949264551173, 
    0.0507689872336721, -0.227836805999881, -0.0274776290627502, 
    0.071949654960056, 0.0963541624731533, 0.396683866573917, 
    0.113075326251613, -0.0445270104397283, -0.112581969403505, 
    0.34694642766221, 0.254325580511115, 0.073422379548652, 
    -0.0676552317639726, -0.0813632219896272, -0.0154501482236389, 
    0.704968330123891, 0.200925093988109, -0.0769909014369915, 
    -0.10888947723161, 0.697342550328149, 0.222038255371446, 
    0.0358516449305368, -0.131501566302314, -0.127993879660176, 
    0.0987082005129911, -0.106759516459831, 0.0817967741406355, 
    -0.111583875586493, -0.00388212861689099, -0.0379203543898036, 
    0.0507963787010775, -0.161892167929136, 0.00217567100687174, 
    0.128362081954001, 0.13516758511704, 0.172016271135027, 
    0.241783634045462, 0.218379950785102, 0.185643688616522, 
    0.215110771759314, 0.203548710034952, 0.200998066307816, 
    0.340828868034327, 0.290280923035949, 0.123680577626112, 
    0.174455955729501, 0.510291456971466, 0.338702233593886, 
    0.0921039543762624, 0.0322201133806849, 0.597460379567636, 
    0.238424900613626, 0.0324480309844154, -0.0829735223056409, 
    0.704035657833186, 0.228724143492152, 0.0168834638827365, 
    -0.133703275767507, 0.0368499424402241, 0.737238862711601, 
    0.323957662608413, -0.0286065410623509, 0.113793232802099, 
    0.361696158613292, 0.408745789336314, 0.23027917858651, 
    -0.0784244050072623, 0.251710876987636, 0.408270192822502, 
    0.399189775184707, 0.00453844726962038, -0.208700165901529,
  -0.0460115427184059, 0.321048625563427, -0.0256208025536424, 
    0.239866335462399, -0.216092848199881, 0.187171196627659, 
    -0.25358396832911, 0.0719814174740419, -0.417171138094336, 
    -0.15984699795401, 0.000556277535472528, -0.0202011496907718, 
    0.0787819369107217, 0.0645565224396655, 0.112942077224701, 
    0.0577690954373646, 0.0693527898490195, 0.124367035436226, 
    0.0805420074507348, -0.00825601966027003, 0.005291999244688, 
    0.131166521739944, 0.251092206027303, 0.186374467100152, 
    0.088300147897874, -0.00180958286158488, 0.121657036533663, 
    0.355993767939351, 0.312888668608708, 0.189837363516487, 
    0.117442067088889, 0.0479430413597773, 0.277759780674865, 
    0.384536498688073, 0.195147952217335, 0.00812797353225353, 
    0.221975969473352, 0.58196824460215, 0.427160605303713, 
    0.198541067615179, 0.0949665903379707, 0.335603531643577, 
    0.461166606218051, 0.268078693576417, 0.111502055208498, 
    0.344870037600204, 0.511864477204223, 0.185747486181539, 
    -0.0491775455555535, 0.0265557086898531, 0.558670670511836, 
    0.245018957015305, 0.0312019604240714, 0.551098283769266, 
    0.238195177408232, -0.0674437872993532, 0.0325087867533761, 
    0.637455759904313, 0.059454347436213, -0.099502244636184, 
    0.137751121716991, 0.36682688657965, 0.168053096768165, 
    -0.377153085424438, 0.523079301228246, 0.475189316740694, 
    -0.13910503210022, -0.245329520119324, 0.128906278706257, 
    0.151937525728848, -0.282697762811642, -0.29365936544687, 
    0.111828822371731, -0.176005683168588, -0.14436234068998, 
    -0.00937554408863178, -0.190339642450127, -0.0695375690610139, 
    -0.0319423942285, -0.171312947051884, 0.0900720915645586, 
    -0.314556942505488, 0.0829781069522315, -0.0874246636671214, 
    0.0977597675019101, -0.175647166422719, 0.0613524708088298, 
    -0.0985997845266431, 0.0131872686157987, -0.410464742767177, 
    -0.0552225326626813, 0.0121999582006653, -0.00702066920619519, 
    0.0139474186522965, 0.0909544574785471, 0.0650072243974974, 
    0.0796293847958989, 0.15929649145822, -0.0189150232202736, 
    -0.0733565374461773, -0.235723568273128, 0.625218202564326, 
    0.118710836466995, -0.151392534807081, -0.0189993951859708, 
    0.58839797139329, 0.254099703815667, 0.10614429052795, 
    -0.311644560414206, -0.00887606833778141, 0.722340120879355, 
    0.286201990255299, -0.22838887290916, 0.38529509400874, 
    0.549910917733891, 0.0774381088225267, -0.088452388636315, 
    -0.125996040469209, 0.382970029100928, 0.349188050827264, 
    0.488560459449269, 0.501439337157639, 0.0453622817585046, 
    -0.0792224603918525, 0.134223619673497, 0.254753762566676, 
    -0.061054168355478, -0.0446638124830225, 0.129869556652523, 
    -0.289622422972468, -0.20291594651423, -0.12968569235036, 
    -0.0796772432570654, -0.134980355324971, -0.119754992540708, 
    -0.201310833657703, -0.0774459216002317, -0.136055872791094, 
    -0.0802586139395391, -0.109835403514271, -0.197111031230176, 
    -0.0325143207815285, -0.138822623421436, -0.0203254626326089, 
    -0.237954797543822, -0.0687163033229622, -0.0263471234373108, 
    -0.0316201794738806, 0.138935702875168, -0.257582636911134, 
    -0.0358125388311407, -0.00914275431849196, 0.0126522458354786, 
    -0.00969267708912894, 0.00237202801005451, 0.0871388748059632, 
    -0.0109388371202167, -0.027348243754009, 0.0926628122248295, 
    -0.391550781147564, 0.0341325509320221, 0.419716932511335, 
    0.312749249276479, 0.303221834365291, 0.433172753043537, 
    0.201532603754659, -0.00154524117299749, 1.0646776020533, 
    0.26076758973369, 0.105083150733973, -0.235605474397672, 
    0.261710162673808, 0.487207117971322, 0.845511999221517, 
    0.416807490356712, -0.263245730652633, 0.455351912910341, 
    0.402826619319345, 0.131511107194595, 0.275019481958345, 
    0.42072923821203, 0.108555133055619, -0.0507641659124917, 
    0.144021801821302, 0.246058513156745, 0.0583783815746178, 
    0.0927569869154543, 0.348886529113536, 0.00937558040565462, 
    -0.0475574545021974, 0.0910876139695462, 0.00182096478603132, 
    -0.168735533164585, 0.27184440129698, 0.913395629482111, 
    0.217921013339762, -0.231299494784982, 0.408911156274629, 
    0.386036451435416, -0.142205253095059, 0.011254765247394, 
    0.0892491572394231, -0.624526144471947, 0.534639038058237, 
    0.329857008033014, -0.246184673026195, 0.508900375154348, 
    0.473405298984231, 0.0613445349507715, 0.255864947011461, 
    -0.201501746169724, 0.225718046970032, -0.210465781098991, 
    0.114796007893938, -0.241158773811785, 0.0647871897689069, 
    -0.432537775890883, -0.122378269229524, -0.110126075677444, 
    -0.297247571909122, 0.0989963673729783, 0.0271044864367267, 
    0.0718666882500057, 0.299815920544189, 0.275714928531065, 
    0.184593909756828, 0.243242735076133, 0.304305786669273, 
    0.26819827229697, 0.257628667344209, 0.285826457844678, 
    0.294513844815882, 0.275529805318976, 0.249762690099385, 
    0.246188061324146, 0.254256182220332, 0.209409438194666, 
    0.161582975671691, 0.271792590094238, 0.333160271512089, 
    0.193373066970789, 0.125538113162569, 0.10692124610146, 
    0.122895777078356, 0.133133289011255, 0.10010162652754, 
    0.0567943214003192, 0.0784406000236171, 0.229483041846022, 
    0.117209358999785, -0.00295110456359642, 0.0326933351650981, 
    0.0905940132620152, 0.304111053526768, 0.494377759726638, 
    0.200497058513903, 0.00767611709051062, 0.0785848989839971, 
    -0.0920341280558265, 0.221685072171482, 0.78480962533444, 
    0.331900624490887, 0.11406786315123, 0.581774140638211, 
    0.213870237533296, -0.375443668701074, 0.310391954461399, 
    0.626395998203151, -0.408959748941626, -0.190069305821184, 
    0.126873670466445, -0.00184660728570565, 0.433872083932234, 
    -0.519065258885359, 0.18555327297395, -0.581147692704736, 
    -0.113888828432609, -0.350323450393078, -0.0632524479936162, 
    -0.35185366036314, 0.0454440206308804, 0.0792060752622074, 
    -0.0758163659201069, 0.0223889201820606, 0.16316998237472, 
    0.0256369379362514, 0.138537529989861, 0.157874711145731, 
    0.0954463370227642, -0.0217015960094388, 0.0432020314619199, 
    0.0896296467709246, 0.136040690008522, 0.121321907730865, 
    0.114577755315746, 0.205436774053633, 0.216044192719957, 
    0.145762838031004, 0.135749488055287, 0.212036379856694, 
    0.241520880069164, 0.202562474397076, 0.183679624490938, 
    0.205996630136583, 0.193264198692042, 0.117816742303851, 
    0.167691729364441, 0.366511924525891, 0.150646665226611, 
    -0.072967641752229, -0.0329968672290265, 0.417368103616679, 
    0.318651063996362, 0.148696550282949, 0.0778179315447422, 
    0.125109597003673, 0.0137927195581299, 0.043307061655998, 
    0.650317656461318, 0.426889050048535, 0.0182522189550829, 
    -0.0377642810805871, -0.268324919185513, 0.328744664000648, 
    0.387035137299136, 0.120988599738212, 0.0191729688145708, 
    -0.175660966464406, 0.33225789319067, 0.345314434593105, 
    0.107033091765359, -0.0165954426997685, 0.298202246965011, 
    0.457962885594243, 0.17931643999355, -0.0303059477980649, 
    -0.0568585747129248, 0.581614452074202, 0.409496892461405, 
    0.0144452274383081, -0.0298307512692946, -0.26293399502968, 
    0.462152145584784, 0.313463183810277, 0.159485228435239, 
    0.165672419781227, -0.110539393616628, 0.593970899382395, 
    0.342909771208676, 0.00844166232516774, -0.348327926800185, 
    -0.00204558546955579, 0.570595587282108, 0.361038360650202, 
    0.132843368808821, 0.110525612165542, 0.538877777063058, 
    0.347204304729786, 0.1309077401079, 0.250938021217063,
  -0.00797483877745407, 0.213301877375602, 0.369391054036372, 
    0.252178191334574, 0.483643658690643, 0.602899725657323, 
    0.242184795757169, 0.0884067594604843, 0.797915604908739, 
    0.468855429652028, 0.0835792513658842, -0.0793112405648745, 
    0.751425492290359, 0.323670123463579, 0.0503937559634231, 
    0.0113969371974305, 0.624521427198335, 0.330448986336784, 
    0.198938307502149, -0.103070062254043, 0.5246461459553, 
    0.430985104852134, 0.272249045831037, 0.0492048865367768, 
    -0.269949677993365, -0.232129518668276, 0.343586837827298, 
    0.398675509833212, 0.593807239812636, 0.41614119193309, 
    0.0667629328719264, 0.465478398136121, 0.0211121180941669, 
    0.0521938091705861, -0.472727608747652, 0.378833333548792, 
    0.387778954121196, 0.133948335693719, 0.00657264733139684, 
    0.265799537540094, -0.249920449608662, -0.2507237814301, 
    -0.269472250982314, -0.105403877764251, -0.281029381631971, 
    -0.0555377330285002, -0.323323423270888, -0.133272359235232, 
    -0.213110096199756, -0.27575891600447, -0.0442869725770449, 
    0.0163106814542309, -0.0068387404659246, 0.00522979621570387, 
    0.0150179552025135, 0.0553182248526555, -0.0320918734129428, 
    0.0370923678241664, 0.0526286167460962, 0.0114181872110925, 
    0.122104825253292, 0.0755679828870267, -0.26219928020188, 
    0.180664760447008, 0.671928939858341, -0.117274746252665, 
    -0.145331856005333, -0.289794405047876, 0.588411614895367, 
    0.28033896521487, 0.0610602290559339, 0.0565026177351824, 
    0.0630897520154564, -0.19820751197355, 0.3999460888778, 
    0.210582626453079, -0.00743080906974965, 0.281919684620855, 
    0.273801728990466, -0.0115449244683179, -0.0744292203156325, 
    -0.124322638248249, 0.0588471835090101, -0.18637288521541, 
    -0.00445490336521266, -0.220407953133248, -0.102703971426913, 
    -0.0530084123567, -0.131551244152867, -0.0257180896361157, 
    0.0343228823524654, -0.0706457047568223, 0.0875741994796249, 
    0.272581650382715, 0.182081523543246, 0.194516828364536, 
    0.254845946143938, -0.0464314465938597, 0.383849645189132, 
    0.406231039693715, 0.460131545119554, 0.265045610477816, 
    -0.00748662210802614, -0.405773914751974, 1.10352742920046, 
    0.622642209775117, 0.255808296536816, -0.180328748027859, 
    0.565457194222589, 0.0730482861394397, -0.419234929924887, 
    -0.0567662001663494, -0.0773813530266787, 0.237359383877371, 
    0.0133697398710253, -0.0529063707330547, -0.0832628446165426, 
    0.057606377487467, 0.286244434802477, 0.191262293986188, 
    -0.00749318545271359, -0.0534514035879984, -0.073434602237454, 
    0.0123291604437695, 0.194566737914014, 0.0735410984169944, 
    -0.0216112221831335, 0.0739358360555486, 0.0851998209185103, 
    0.0231957679541902, 0.0194732903662477, 0.0359218509245306, 
    0.00150318540547273, -0.00321293163932015, -0.00370606628091871, 
    -0.0194214219951616, 0.000822022420759072, -0.0268705783135334, 
    0.00248533565783299, -0.0100942367341197, -0.100847280554571, 
    0.00996401788316569, -0.067414189303932, 0.0354096152118048, 
    -0.144067100593822, -0.00748011946771333, -0.0982903540448195, 
    -0.105047071187879, 0.0544903936946612, -0.112730797707161, 
    -0.00475010679922114, 0.0634166172275446, 0.0986286447063168, 
    0.101263035684764, 0.108272416712525, 0.10383040757845, 0.15918378144078, 
    0.29610234657085, 0.200071036711594, -0.225966932652417, 
    0.415544342760627, 0.366547822612741, -0.0173059021670553, 
    0.342445141621506, 0.489012790705853, 0.108343591263794, 
    -0.00294150362640987, 0.541255302236874, 0.647260702231926, 
    0.224838903750646, -0.00276140975628483, -0.18257572070851, 
    0.303597582645719, 0.368853691660189, 0.311076827751839, 
    0.379124300172628, 0.201406286678446, 0.258009531664873, 
    0.766733840805425, 0.0274039362310035, -0.119230380389371, 
    -0.0133589609413771, -0.0841530928912219, 0.0712742527113157, 
    0.113439162478742, -0.0939428635589358, -0.15874082991168, 
    0.0335500463531819, -0.030108306810234, -0.143106473892382, 
    0.0470060229273314, -0.111702297647783, 0.0390855668357221, 
    -0.104264896290731, -0.010131574032574, -0.109286669950198, 
    -0.0884015756098414, 0.037381255427623, 0.0507636218404885, 
    -0.177427922966826, -0.0437312586226186, 0.274880391911248, 
    0.0371121685143908, -0.031882119067016, -0.126134471227081, 
    0.328082086267233, 0.25515581695318, 0.0344269927049239, 
    0.0421606360250203, -0.0597504005695653, 0.714156726826388, 
    -0.0855036119260232, -0.115533011034882, 0.081414120305239, 
    0.128595449057121, -0.0488071921301365, 0.685242303995637, 
    0.302074513105539, 0.705950724850114, 1.19955295741809, 
    0.0491044389848631, -0.153798720745458, -0.198116149223379, 
    -0.102694030407476, 0.234626847116685, 0.135746372207279, 
    0.0645352882719332, -0.096947688556848, 0.170537165853889, 
    -0.0430447055190633, -0.156373237528539, -0.0598208746740879, 
    -0.0985074042727476, 0.0247073972910614, -0.0760668994840839, 
    -0.0193004968467948, -0.0347065052760823, -0.167590457860715, 
    -0.0194394473134091, -0.0764872475557736, 0.0810150512861062, 
    -0.116268013112355, 0.0406113434822827, -0.0374078300098329, 
    0.05233932327845, -0.105046222148397, 0.0345399211946979, 
    -0.00597401583104201, 0.0814852760368977, -0.186406700262967, 
    0.0602479237958804, 0.0954778590955892, -0.0208297055911306, 
    0.090035703408774, 0.282752549322302, 0.14887906177925, 
    0.0555239154453813, 0.0791503968196187, -0.205095706573144, 
    0.445896574251674, 0.326210367876188, -0.131090512841872, 
    0.405046088295521, 0.548102549552238, 0.10523215907964, 
    0.310332562673964, -0.318674487785055, 0.111647126997814, 
    0.600214295979473, 0.133679881645074, -0.057894532755596, 
    -0.206131955409642, 0.502171835099523, 0.292984331611785, 
    0.118789176565298, -0.120342913964572, 0.21850135732643, 
    0.16471196942536, 0.505702621662884, 0.579571153931289, 
    0.054353540147082, 0.0116871091911244, 0.237048171865974, 
    -0.158547450368237, 0.0132925721259916, 0.303593749061544, 
    0.0452565316779374, -0.112766824959112, 0.0288527015280338, 
    0.295983948568996, -0.0494036523274325, -0.00271335497220432, 
    -0.0287251959736591, 0.00171910602004023, -0.03257223306341, 
    -0.00457385954628628, -0.0410743834973854, -0.00297911247169046, 
    0.0915337038356619, -0.130710229267833, 0.0906161479001609, 
    0.256598815645472, 0.130320018181436, 0.0581562876265129, 
    0.0421623959629811, -0.00995151761750414, 0.436061596394261, 
    0.663853851149513, 0.0526343011522414, -0.364874686227719, 
    0.0287896473261945, 0.562784612726441, 0.179394160410992, 
    -0.228843970415403, 0.419808384143811, 0.749597116387056, 
    0.323272512139718, -0.0272169394707465, 0.697267776407951, 
    0.433588710435577, 0.00627529654310743, -0.000407811033052832, 
    -0.205468694144666, 0.34927418456358, 0.224573752769142, 
    0.137593878701689, 0.154532820304231, -0.00505136476255792, 
    0.470262533445101, 0.00283320697569124, -0.107817561606159, 
    -0.225187313622915, -0.0207258355936988, 0.0361021994245817, 
    -0.0922540342927651, -0.0653229800302361, 0.117940166470152, 
    -0.127879711447784, 0.0505548444896134, 0.056661877417519, 
    -0.0535096886180182, -0.0137512285182163, -0.277072421654044, 
    -0.0389954628607071, 0.0282364786966577, -0.243978660868854, 
    0.184041800345525, -0.0539672405358243, 0.0505433720617825, 
    -0.237647133020378, -0.0111162113942961, 0.0742689360766067, 
    0.139325711263485, 0.132148227533484, 0.102332326245218, 
    0.0973968519978538, 0.262421172229157, 0.384279671711799, 
    0.234392699949867, 0.0777632308714986,
  -0.00563792712966432, 0.564379639748641, -0.0351843165143208, 
    0.168906321335061, -0.352171874230875, 0.498925456735744, 
    0.233897384513467, 0.127286708090979, 0.305615111437527, 
    0.231350341080405, 0.0535976269003413, -0.170630059258302, 
    -0.117945475097687, -0.0953398816365155, -0.115237926014925, 
    -0.0614111216164157, -0.0978277698465401, -0.107809865191203, 
    -0.0736401200740809, -0.131251088422388, -0.00999941484458269, 
    -0.00278057437582599, 0.184049183149925, 0.228147340807198, 
    0.121316330286727, 0.0224767840511441, 0.102601944223052, 
    0.288890514254246, 0.143005017252799, 0.0173397949319795, 
    -0.0110188220690355, 0.327904289258819, 0.21835996997421, 
    0.0351098091083862, 0.163755394531469, 0.343995363925698, 
    0.167560663593121, 0.0459549467342777, 0.33528378006029, 
    0.316661453978508, 0.113660060547211, 0.0723405957375536, 
    0.0817902628473572, 0.0879448375595274, 0.0942893513846331, 
    0.104884903963347, 0.116532761876802, 0.0983668824460948, 
    0.0746535259812821, 0.0151503630400859, 0.2676436947509, 
    0.183203496431596, 0.00953641732317946, 0.333687001091522, 
    0.320083791433849, 0.112482835322905, 0.01669636407287, 
    0.433901976022695, 0.241877363059509, -0.198139241773131, 
    0.353218970974606, 0.553635470880502, 0.209454019261579, 
    0.104572865636825, 0.161526967737074, -0.29808075948961, 
    0.339870499926717, 1.13012358244358, -0.180062818696476, 
    -0.115150646077976, -0.197284415089213, -0.249079890181201, 
    -0.144014128206324, -0.147951821471196, -0.240344379359717, 
    -0.0891541587356241, -0.384832657326774, -0.149633882440565, 
    -0.167826443520256, -0.227048281998647, 0.0434064478813922, 
    -0.114474507858237, 0.0219890685764756, -0.0436392172978653, 
    0.181589145521189, 0.114928362618713, -0.0395913758196646, 
    0.119393303477106, -0.271480706631306, -0.0511019593183112, 
    -0.0386201222963829, 0.0286264259407026, 0.00520274146582199, 
    0.00900371588460072, 0.0191407967178843, 0.0359209558665349, 
    0.0252080011622978, 0.0160331971990734, -0.0306988051233504, 
    -0.0324583450190887, 0.0495303478807751, 0.0944786015577806, 
    0.11105171810207, 0.139486441237994, 0.149229235569063, 
    0.0879246396159155, 0.0855492375130593, 0.277995326814926, 
    0.0964413964221713, -0.124188268632342, 0.0319326560682367, 
    0.460004476412484, 0.0835299379893835, -0.0923135643688764, 
    -0.104915628911876, 0.288574475306833, 0.535379889770629, 
    0.271780244919636, 0.102234709434586, 0.495213245822958, 
    0.161953821729646, -0.0558806461641035, 0.181394188808497, 
    0.353165590019939, -0.184739670373076, -0.236461731946502, 
    -0.0714038644959996, 0.337388672666497, 0.0729644366589218, 
    0.0183694865640072, -0.0400193903397402, -0.302190627299507, 
    0.0589631461435273, -0.119231252521426, 0.0164409273236739, 
    -0.226229015096996, 0.0196077146294058, -0.179048120353262, 
    0.023178673855108, -0.294227976198895, -0.0235826113030616, 
    0.0522875434367593, 0.0871500785283752, 0.157359437157929, 
    0.224518945011046, 0.157650322350174, 0.0880969526324907, 
    0.210610751393183, 0.244803370844509, 0.127626476305923, 
    0.0885884043439196, -0.0660996330868588, 0.33997704414065, 
    0.531618167419471, 0.202081753798826, -0.0316209700208511, 
    0.165984351626872, 0.356777992293746, 0.113253391400392, 
    0.570609506288589, 0.626567867473012, -0.00173907190224343, 
    -0.325619726516602, -0.0101306994342775, 0.9746163571698, 
    -0.00563845221974571, -0.0438719667221623, -0.0611629423297293, 
    0.634309766898853, 0.0833332315196488, -0.0231713737491447, 
    -0.216592208581572, 0.0701231491070532, 0.225406964907032, 
    0.065621229741268, 0.387858809355822, 0.330735228054232, 
    0.0668127120195246, 0.435136088514894, 0.109337667434321, 
    -0.234580666411402, -0.01125717331379, -0.140307488298868, 
    0.0119938013452826, -0.175839292852721, -0.0504095805810764, 
    -0.11201883529553, -0.0980438345124248, -0.169085968385398, 
    -0.00374831611384307, -0.0953091307808367, 0.119097095086831, 
    -0.0359560515075734, 0.0610093674407613, -0.0734261596155188, 
    0.0385471311682188, -0.0611916501714435, 0.0150597165185558, 
    -0.134210702779968, -0.0446862164814418, 0.0157284179616876, 
    -0.0623308202473443, 0.0184416230148652, -0.0288986624681246, 
    -0.000420623477202925, -0.0433972208376472, -0.0235408055161099, 
    0.0214424652807801, 0.0760869698964881, -0.0868608669599293, 
    0.0728454727756525, 0.161415463855075, 0.0724291740010066, 
    -0.008012392141435, 0.115437255962312, 0.239007076998816, 
    0.171410861803858, 0.139136947899457, 0.221283733593185, 
    -0.316026342141167, 0.53108538122238, 0.355828298620073, 
    -0.330757710866984, 0.587495339701949, 0.490126087907698, 
    -0.345514513105521, -0.0314236260539562, -0.196229405266407, 
    0.838218473858068, -0.136306814024031, -0.190599080024757, 
    0.0173185177698747, 0.333244348148218, 0.000367287623859777, 
    -0.0138336938637013, -0.106082300141438, -0.06645947887495, 
    0.523650570634246, -0.0276636380696804, -0.350010156604016, 
    -0.330461401593818, -0.136119598393814, -0.150591380472712, 
    -0.0675585483189277, -0.289888553497058, -0.0241228751939636, 
    -0.279815214862933, -0.0580528269758691, -0.218432005724623, 
    0.0205481829101139, -0.119934446555534, -0.0167525098867877, 
    -0.101882981059662, -0.195231401647572, 0.0862185114291849, 
    0.00932956170985733, 0.113321807328469, 0.0174661643548837, 
    0.0783691527075776, -0.118517352226191, 0.0103042815072699, 
    0.0117374944158511, 0.033112039118843, 0.0120789326796704, 
    0.0248749528571148, 0.0139209887695606, -0.0163071973343352, 
    0.0973048994902145, 0.0970367001553564, -0.13615458259242, 
    -0.0681396044323306, 0.242712372840283, 0.362877264000938, 
    0.209932680162306, 0.0387047973284459, -0.195763441050265, 
    -0.0523096395513139, 0.599385371431414, 0.0722555679778353, 
    -0.122761743588665, -0.00158945302512183, 0.106654279425014, 
    0.358079874531064, 0.69692280522285, 0.522339912271131, 
    0.212728131480142, -0.41222312439378, 0.390353693610478, 
    0.495476112254532, 0.209948103744298, 0.164261932269798, 
    0.42722680152289, 0.143433268496687, 0.120776643370004, 
    0.139332494769738, -0.16453079858034, 0.311639340357834, 
    0.219408653909263, 0.0452414321575106, 0.247361908204863, 
    0.215386970841111, -0.0132141978894535, 0.180295828962409, 
    0.327752501386421, -0.0105188304444661, -0.0306446128264623, 
    -0.11632250205865, 0.228818533908092, 0.199965060866042, 
    0.0857035413819602, 0.0631824031831962, 0.165636090110204, 
    0.0149161991750143, 0.0233285939515768, 0.0525497254639456, 
    -0.065162942526048, 0.0652700942165282, 0.121478326482335, 
    -0.0483203923521998, -0.0468750073472236, -0.082488539286531, 
    -0.134982353148317, -0.0453173842658117, -0.0288620724747139, 
    0.0467569189463014, -0.0489009821906547, 0.103970203443949, 
    -0.0705385137353801, 0.0945391692880765, -0.169921531995889, 
    0.0791022850779274, -0.00655026288979459, 0.173133319116595, 
    0.243840574199882, 0.0835549593067923, -0.0964129127118954, 
    0.0615586175836736, 0.3922685139647, 0.116192420826985, 
    -0.0043516912962035, -0.0157924180755566, 0.654342186599264, 
    0.0484174995691343, -0.0880306186516015, -0.281265767721616, 
    0.777747015705204, 0.232187150707646, -0.192955410153792, 
    0.361296978567054, 0.584743785996387, 0.196305595996638, 
    -0.110897837570737, 0.596154949504527, 0.611364815846812, 
    0.0513285767107229, -0.457357262175262, -0.0399403937991013, 
    0.63672047862208, 0.161761705032265, 0.142252360665883,
  0.176665532328233, 0.105805264836527, -0.0257277918385331, 
    -0.298655181617542, 0.391346745541432, 0.256201316815438, 
    0.0707757237682339, -0.191285409944464, 0.153878481922663, 
    0.379177200350436, -0.0206421828503502, -0.0259283439157936, 
    -0.090943136004915, -0.0557217975009493, 0.287893576285595, 
    0.202926646425622, 0.0632022923929788, 0.204133917986893, 
    0.0705893331210348, 0.226037353816791, 0.482895374139667, 
    -0.0497698866399394, -0.071752521151375, -0.338759173953798, 
    0.178189999243103, 0.572024922740581, 0.21214128327006, 
    -0.149135490382561, 0.179242860164881, 0.419441373837862, 
    0.110715397585341, 0.0408132322231832, -0.0246817263747201, 
    0.181321155064014, 0.309727250994619, 0.204398676757564, 
    0.101768613722693, 0.0656109551000849, 0.224352076676857, 
    0.260523029559819, 0.116714330913609, 0.0604691797597282, 
    0.443243873409394, 0.304705124917772, -0.00282764289574067, 
    -0.124659460199854, -0.164677061101242, 0.348983240379074, 
    0.245359448225889, 0.0998788345375481, -0.0491871843459833, 
    0.175502816798472, 0.154050199227621, 0.0864954957314999, 
    0.0856839468012342, -0.0010266914179913, 0.115582555933677, 
    0.313829210336493, 0.114971094210081, 0.0190731336815557, 
    -0.123486584846614, 0.0437743280787854, -0.112692427966699, 
    -0.0141544387802847, -0.0352688122518423, 0.0291285953064611, 
    -0.173956509870693, -0.00997116526402006, -0.14861135306859, 
    -0.157493955911498, 0.0147351670400831, 0.106062868619909, 
    0.0690657533652705, 0.111576467474165, 0.263589999896525, 
    0.155808988179595, -0.0283730481029412, 0.242759722963229, 
    0.326608394067087, 0.160198122778385, 0.184114488936087, 
    -0.281775446726372, 0.107507084183859, 0.60010281953829, 
    0.115226269111825, -0.0146231381853758, -0.239727082975599, 
    0.23948697957082, 0.469110842211544, 0.463187403008389, 
    0.153621727443814, -0.328362003480901, 0.137685584047359, 
    0.227378305199074, 0.216784675903648, 0.606846620371055, 
    0.161172387689646, -0.12524292001562, 0.302005947224565, 
    0.256609455965123, -0.279148697590312, -0.140266873875486, 
    -0.0581817040170673, -0.152516013546068, 0.0592925173651955, 
    -0.307873631784995, 0.044337467517341, -0.478878867696287, 
    -0.251931438957738, -0.123058463653618, -0.408287854386196, 
    -0.0161257767138952, -0.164670436116409, 0.0504080683199069, 
    0.0370679023098864, -0.542660034159163, 0.0330181431407705, 
    -0.0508523488054567, 0.0960056762594978, -0.331459762704593, 
    0.0174812088645967, -0.0111786642545666, -0.0126188093571129, 
    0.00335925538197293, 0.00531975611846533, -0.0174047778661595, 
    -0.00985318985405499, 0.03654836230288, 0.0260291835037181, 
    -0.0638842728002896, 0.169560112675925, 0.13474289520212, 
    -0.0217735829417817, 0.148922077508195, 0.39542726971352, 
    0.199814870758988, 0.0541770452241674, -0.0755695385881832, 
    0.148958335049803, 0.458418387493043, 0.264699275257182, 
    -0.0872795114833791, 0.328937480725152, 0.453249768180481, 
    0.0412849853629412, 0.285438457411801, 0.62137893723602, 
    0.518162221529996, 0.376547275712742, -0.0243222731781844, 
    0.675039004743028, 0.236380855124552, 0.0268655791821889, 
    -0.199877280783496, -0.0581567494489616, 0.767144259045324, 
    0.174234206538136, 0.0119299584352554, -0.220293469943641, 
    0.424008787081562, 0.417512040695084, 0.0409775198679947, 
    -0.0777965088093616, 0.138932468210908, -0.191400230795535, 
    0.55693866950916, 0.239302032247214, 0.0206887053417883, 
    0.354001556887678, 0.141455111103314, -0.161105516543184, 
    -0.147165800763575, 0.0199517014025279, 0.058103885716464, 
    -0.0128943799601351, 0.00594700043869606, -0.0785120624062126, 
    0.0105924443444409, 0.0351862916569059, 0.00736689280502401, 
    0.112153971997982, 0.0745245469755041, -0.0232732112056605, 
    0.13142852838919, 0.271968480421059, 0.145375826147933, 
    0.049034020188879, 0.0173800853514578, 0.0965123514666303, 
    0.33275609663505, 0.288017425986725, -0.0106528073935121, 
    0.212354297452101, 0.52759099933694, 0.101233229204963, 
    -0.356362400120313, 0.376404946865517, 0.76939163896235, 
    0.192973795874947, -0.121577782338356, 0.0127419537560396, 
    0.336502796422358, 0.435893636443915, 0.199471535262534, 
    0.349021759787198, 0.772759523825575, 0.311131681715587, 
    0.18568036170063, -0.150082694498726, 0.415394216758473, 0.2946168358645, 
    0.122168701911694, 0.0759136425436328, 0.0766812026818662, 
    0.0744763456409082, 0.0613831135669556, 0.0246916303310751, 
    0.159028971681224, 0.0687128406599472, -0.00704577864371617, 
    -0.167625069828506, -0.0139576174964848, 0.498791499064455, 
    0.205710174068048, 0.111369404378593, -0.148169469044058, 
    0.279272939995621, 0.353253205336594, 0.396090511880506, 
    0.218229841078758, -0.137569500663867, 0.198900687683466, 
    0.333957898894907, 0.346001388233853, 1.2551325229492, 
    0.0593894967069922, -0.239604820478714, -0.0446488376051621, 
    0.938156393880671, 0.0639238708310362, -0.162538538537223, 
    -0.126774239872451, -0.0204572935719086, -0.455183699138582, 
    -0.153033522063046, -0.21364314632171, -0.294235736982244, 
    -0.082409720073921, -0.320297466691043, 0.0811368200407146, 
    -0.114303533173445, 0.0919797345778451, 0.0853267901835721, 
    0.137611939972588, -0.196180138005985, 0.0440310374011391, 
    -0.0986981295491865, -0.15916646493072, 0.0775507908693499, 
    0.0247305922668419, 0.100634825160323, -0.102013264383013, 
    0.0254256736075076, -0.157898184442522, -0.0167225228492814, 
    -0.123482216102871, -0.0117040030697946, -0.119612333398219, 
    0.0186536881204752, -0.206024095210969, -0.0178701793260009, 
    0.0217279394343168, 0.0405076837721903, 0.0632751014285092, 
    0.0790644376510334, 0.0592282822539598, 0.0513377447506695, 
    0.110311989486591, 0.0962971182244257, 0.100723264268412, 
    0.203825156136726, -0.0227868869369235, 0.441996521604778, 
    0.244115519108963, 0.0613622249745275, -0.104708268514391, 
    0.427734155426169, 0.303021523267482, 0.107358389769445, 
    0.0170374067356223, 0.103928223964009, 0.284009618172406, 
    0.30888585252685, 0.286414168585726, 0.267047580718109, 
    0.225297028363951, 0.217463454016389, 0.249895679150366, 
    0.206324588673916, 0.154473560831331, 0.283665927138484, 
    0.341004423049399, 0.184245807874844, 0.024785061158439, 
    0.111061497335187, 0.408948468553765, 0.374434964545402, 
    0.283401882239007, 0.161255824721227, -0.129963454323081, 
    0.247843005876186, -0.0509542437837242, 0.371916156046099, 
    0.991200314182704, 0.0425986995229413, -0.165242887299867, 
    -0.0351283226033061, -0.112819087004109, 0.78378153639618, 
    0.664257837774313, -0.0262829446420878, -0.117389770490558, 
    -0.0877299740571005, -0.0888713498616301, -0.0722585088677378, 
    -0.0797449561893115, -0.0549016741246474, -0.107511614609271, 
    -0.113569157239927, -0.0467506527820192, -0.0543025941068032, 
    0.0371915828626784, -0.0199927082272656, -0.0269962847432377, 
    0.0706322630325376, -0.0264092187947673, 0.037102333940046, 
    -0.0104988325205433, 0.0358294578915277, -0.0563053130350539, 
    0.043239439639458, 0.2139646680736, 0.231497400968127, 0.113684788433866, 
    -0.0362096236779385, 0.0804349791666077, 0.193500082768193, 
    0.174963156689369, 0.327573333359333, 0.434390382066846, 
    0.40398983609264, 0.223619458494705, 0.122693081905298, 
    -0.105199487301677, 0.294057258712383, 1.12397878972283, 
    -0.262282268973461, -0.152663924202363, -0.0865743897555469, 
    0.895493719947363,
  -0.059674166385206, 0.0968840570064023, 0.128209706658137, 
    0.120858758016977, 0.158797609973029, 0.150090637616483, 
    0.235916072780027, 0.387546554452218, 0.191342080990778, 
    -0.0611683222335797, 0.0186170773008147, 0.670974899397146, 
    0.294338217150829, 0.0573562043737991, -0.181083075232521, 
    0.620949314373679, 0.461441121740361, 0.184544303089751, 
    -0.24966586256962, 0.463768161506975, 0.524780122866028, 
    0.0977900245191947, -0.298024951569698, 0.0996766336562369, 
    0.508058149395917, 0.101235084069257, 0.0962186100058612, 
    -0.247751339741382, 0.342267105360784, 0.33522580322973, 
    0.0287461086070025, -0.0347135637655502, -0.143265493515449, 
    0.0556586079213326, 0.213053014244452, 0.533827591485271, 
    0.208129093541138, -0.13571838517239, 0.233211680384722, 
    0.284113541879364, -0.168634553188574, -0.0501376207482235, 
    -0.100469799316815, 0.128413434452061, 0.198921818408329, 
    0.118074568548203, -0.113176956273286, 0.0218701508114457, 
    0.179239674847045, 0.0385455111928761, -0.0315447606224274, 
    0.139517875123403, -0.0674299892626209, 0.125598661985348, 
    -0.344691264766961, -0.00771369823708863, -0.215379798323315, 
    -0.175755400219003, -0.0381286047202254, -0.174153101465698, 
    -0.0173223817820152, 0.087211842221005, 0.0527935128392611, 
    0.0687298519711662, 0.101408026160833, 0.0620344376301574, 
    0.0718297755658092, 0.109339333038194, 0.0951387608995386, 
    0.0354013920031611, 0.107124172373101, 0.162136758026823, 
    0.166327048766029, 0.17881060626681, 0.174535992530484, 
    0.142659164146647, 0.295102914439582, 0.356883387273468, 
    0.096994288947912, -0.0590710916045115, -0.169357398411942, 
    0.41184278723191, 0.43890281104109, 0.189095284250921, 0.182276957883504, 
    0.615016394851596, 0.104756512534396, 0.0892371635487691, 
    -0.296050629487546, 0.196283628149633, 0.417818834998429, 
    0.272802568697422, 0.11569888052195, -0.024332214806029, 
    -0.192522982589022, -0.0660277566655248, 0.370698869133205, 
    -0.0865692471163439, -0.0305924744473498, -0.0478281376472735, 
    -0.170240405069807, -0.24305176850644, 0.118921915307016, 
    -0.146948398981076, 0.118599726434497, -0.164198410592792, 
    0.0564902467447857, -0.110852359871916, 0.0519132892974907, 
    -0.259352408677981, -0.0112296868296588, 0.0535498642853461, 
    0.090722714622486, 0.144751749355262, 0.151356264286661, 
    0.102599137967218, 0.0943282070013458, 0.148511260851641, 
    0.128169038243051, 0.0468495457273599, 0.106847635618526, 
    0.226456870341081, 0.183281942879881, 0.170806467709218, 
    0.269192871464689, 0.198965300555972, 0.197044251666166, 
    0.337183322056873, 0.170696191588617, 0.256826032375324, 
    0.62122745290014, 0.0548625950176922, -0.106855427982087, 
    -0.218565255294373, 0.261912311349923, 0.425832352604856, 
    0.226382431584654, 0.342996339415401, 0.749591091122133, 
    -0.139447678025093, -0.254860756894234, -0.0805316597490362, 
    -0.195671238749686, -0.0645582605412379, -0.21905943845817, 
    -0.0476129123287955, -0.234666405603038, -0.133594368422852, 
    -0.0436458271357996, -0.20464996973686, 0.0973530415312991, 
    -0.0243985606752858, 0.028422973254418, 0.0244817506096219, 
    0.057360802558087, 0.0335049507526368, 0.0710024940119093, 
    0.0117647613807054, 0.0345697624661426, -0.0491678066395403, 
    -0.0122444690531228, 0.0685395579891, 0.117655795084475, 
    0.0841344412063321, 0.100099522301943, 0.0997049679140176, 
    0.00500579943873279, 0.402707425750162, 0.268202504297873, 
    -0.159030856095963, 0.438107466449671, 0.291446348143528, 
    0.0712782960266432, -0.436121906487962, 0.303175621096308, 
    0.566993631114972, 0.291295791166646, 0.131097161893129, 
    0.728857121592579, 0.157444382661685, -0.0777731676058557, 
    0.0463860807967973, 0.150283996889553, -0.0269319344609335, 
    -0.0793815323654315, -0.0680628074772571, 0.156676877926402, 
    0.117398358247831, 0.0795971431228618, 0.0750635462592891, 
    -0.048032886383249, 0.08238535516663, -0.00796625847862988, 
    -0.00660793358752319, -0.43878228213124, 0.0314723877580042, 
    -0.235108235061375, -0.287279797852906, 0.115616855651105, 
    -0.283737432644661, -0.0600895311333751, 0.0902537472432358, 
    0.0411382446943837, 0.0819253488304036, 0.0540889283374796, 
    0.0332935557965903, 0.0993697337743058, 0.103357570452681, 
    0.0895935431771972, 0.123757921205311, 0.0363608690467932, 
    0.0494629584929641, 0.0565959022157911, 0.0562277041546542, 
    0.0593401275906527, 0.0495178651242967, 0.0908894060270457, 
    0.0621366175835611, -0.00341559391192028, -0.0213096539768339, 
    0.0322542351835339, 0.728891962346919, 0.219667588825049, 
    0.143223359823136, -0.341708007052641, -0.0160512146116835, 
    0.834345520814072, 0.274981039554416, -0.259102476265058, 
    0.171284564900824, 0.448530727972518, 0.222939261687452, 
    0.112194053403099, -0.169212308356337, 0.090110290401615, 
    -0.133198236388494, 0.614202115064337, 0.486783449548362, 
    -0.189873883524206, 0.014996411186283, -0.309681004894734, 
    0.113384112206226, -0.200106742080774, 0.00834535051173565, 
    -0.3330337284561, -0.109674897888033, -0.139617340502822, 
    -0.232592567529679, 0.0680868326230146, -0.222182999950269, 
    0.105491693124352, 0.0633275324237634, 0.0917146472307133, 
    0.215981710622143, 0.313752273669036, 0.30459451022311, 
    0.176910444677742, 0.0328724649608259, 0.213702127422782, 
    0.379719662010322, 0.240039120526603, 0.165929617621418, 
    0.150441589396991, 0.129787814590873, 0.0851344843690127, 
    0.0940465963461104, 0.0908748928030854, 0.127988858397453, 
    0.148501578531636, 0.0979412291929011, 0.113333905670306, 
    0.103863216748531, 0.107504986701467, 0.238996281563666, 
    0.19952965615629, 0.0297939894404683, 0.185885941968313, 
    0.377539560020371, 0.0170542945180385, -0.0691594765234568, 
    0.0584578767037256, 0.371284855026478, 0.0819731677271769, 
    -0.080899346053175, 0.316606524249309, 0.683513221736808, 
    0.503762571627362, 0.135176506167695, -0.0237603246317062, 
    -0.428490746739053, 0.111390070616879, 0.83474038575765, 
    -0.0123838978262652, -0.144692346332402, -0.170636649159323, 
    -0.133947481442905, 0.0882040555095908, 0.600166076399697, 
    0.107794379911781, 0.0261219605777191, -0.104436089974209, 
    -0.239562374517291, 0.0414769163848084, -0.131131984243525, 
    -0.024862726944426, -0.0761201833664084, 0.0250205765426001, 
    -0.061488317725161, 0.0886067014499917, -0.206788053228063, 
    0.0527345043951308, 0.113446628709678, 0.0903755650957819, 
    0.215405393113448, 0.322503303783542, 0.254634364506539, 
    0.178594357327763, 0.12660804069218, 0.0969943743444695, 
    0.512653956678807, 0.554884518044564, 0.176201404721489, 
    0.0629169417132493, 0.928421482049846, 0.213276381829697, 
    -0.330437917082493, 0.177276210094417, 0.812559997956397, 
    0.157065080338105, 0.136482844758172, -0.27450368730252, 
    0.39041637126459, 0.327650919671833, 0.317293161894025, 
    0.498880226808721, 0.0749485046363496, -0.125795835538722, 
    -0.212002272310871, 0.0384594428292942, 0.614258921230898, 
    0.439364234146792, -0.0260817473788501, -0.20969765126277, 
    -0.195263073944575, 0.439548922864947, 0.187205132004479, 
    -0.0103245039115148, 0.217818979185934, 0.314160199036647, 
    -0.118197740038261, -0.0792249493837104, -0.222990492289423, 
    0.00274758608614561, -0.0790608741740885, 0.0188407473871861, 
    -0.206783126083655, 0.025058479753291, -0.136209083473949, 
    0.00705424749969813, -0.268512951996304,
  0.00539154102896282, 0.0395631988740913, 0.00905987416580092, 
    0.0287419383766908, 0.0091784017918739, 0.0132043407003892, 
    0.0204745068693304, -0.0118829821057743, 0.0766519551120069, 
    0.236945706656793, -0.00691822812640776, 0.022266544251813, 
    0.498338285795375, 0.727836727653722, 0.0837824813284533, 
    -0.185332721883248, -0.0695468155653509, -0.0894278550119015, 
    0.482404868553962, 0.498421739394711, 0.104421792705729, 
    0.416888656242429, 0.535731329349389, 0.0963058872890432, 
    0.0268570510307127, 0.0602690442390227, 0.00403102643655033, 
    -0.226154905866431, 0.149528781662829, 0.233457061320615, 
    -0.00548847520349273, 0.0139144359032735, -0.0654180440735924, 
    0.0292116960249436, -0.370700033070255, -0.0297722313414944, 
    -0.16391124972314, -0.22791997724466, 0.149772229224524, 
    -0.298000198646508, -0.0259848004000038, 0.1313355104924, 
    0.077040919387243, 0.0759681674455597, 0.405625602915739, 
    0.301877247705685, 0.0740961711634149, 0.00823559654301828, 
    0.44336840242861, 0.361243550243336, 0.151095098712736, 
    0.109760250759652, 0.135563500450584, 0.125343140852144, 
    0.126239430921919, 0.110709540644337, 0.114131928384305, 
    0.17191952473636, 0.165474480496634, 0.107135868561216, 
    0.109237284010436, 0.120085415915117, 0.096571074139809, 
    0.119738406865705, 0.192829304006653, 0.177932247198303, 
    0.118805204081936, 0.154043134752815, 0.198068616819239, 
    -0.178771398424096, 0.521227053203044, 0.387584103185398, 
    -0.155942269344469, 0.307228625092657, 0.715210343780752, 
    -0.0810261462752954, -0.130324765173953, -0.184613129281628, 
    0.406371764434738, 0.337780131537854, 0.324701396053804, 
    0.347707694948439, -0.00682894585972069, 0.0313527642929455, 
    0.703034738906253, 0.133939565426981, -0.0600045610675546, 
    0.334118377188632, 0.273726984887876, -0.0118156544016031, 
    -0.319530757456331, 0.0897503896939378, -0.0959565169367395, 
    0.0643342516490692, -0.291970595343588, -0.00649253039469053, 
    -0.591013060545552, -0.24521830621649, -0.0584883059855921, 
    -0.38115514462646, -0.105974088382796, 0.105281840450914, 
    0.106387351137169, 0.149302390878985, 0.102055689672424, 
    0.0330475395627179, 0.0427770688927871, 0.163257085438004, 
    0.148060392115627, 0.0835900547603559, 0.129232278223721, 
    0.132132579532751, 0.0948346952572778, 0.130876529221314, 
    0.272597009483523, 0.169683176084257, -0.0361445115741867, 
    0.226437466713513, 0.274247100615457, -0.00162544539387661, 
    0.292808367060384, 0.346344799677409, 0.20717661572935, 
    0.333650987785396, -0.199767291059307, 0.591748538341513, 
    0.965354159300897, 0.0859350078082776, -0.0294547095360433, 
    -0.0861181605018439, 0.37082603657695, 0.196317309463947, 
    0.0693683507443062, 0.0455474648426946, 0.052472841554033, 
    0.0502350182314977, 0.0518926778637771, 0.060153115381177, 
    0.0516702874630625, 0.046735926405695, 0.051973504341944, 
    0.0451150775707457, 0.060400763762862, 0.0475738431768043, 
    0.0542378254789849, 0.0440909061127078, 0.0515458902683194, 
    0.062793632961528, 0.0614648315513554, 0.0187331606594194, 
    0.0779747317723879, 0.103127408294469, 0.132967500835988, 
    0.160268138577756, 0.131414130309709, 0.0745474370570845, 
    0.131319765854007, 0.250371112398095, 0.174296184367506, 
    0.215337380995152, -0.454233726188417, 0.689205225936474, 
    0.409046013241813, -0.245089359630692, 0.072979166201596, 
    0.861870019916245, 0.270380518829954, -0.00907584298013037, 
    0.328875991918149, 0.456954279851124, 0.195143016711837, 
    0.201502556752582, 0.235898515091532, 0.186307910818829, 
    0.162802584392144, 0.178938495517776, 0.150490588393361, 
    0.104689480995912, 0.165780786353254, 0.229015536914828, 
    0.156961307233915, 0.104451264202589, 0.0800021871700619, 
    0.092791934305302, 0.105211964866738, 0.074823150842428, 
    0.0722814916518286, 0.128771625642805, 0.104778704717648, 
    0.0542368683232081, 0.147368356441494, 0.164727394749029, 
    -0.19802343641663, 0.132753111057054, 0.596902765787623, 
    0.192302636203246, 0.00394279376399996, 0.272653879888137, 
    -0.0232606006392319, 0.38665998748475, 0.768215430831658, 
    0.222843419325618, 0.0175454511688066, 0.31529393953006, 
    0.500320238439956, -0.212523126077921, 0.156364609573202, 
    0.746603954273331, 0.369955971765286, 0.0996337449944375, 
    -0.0994932421655487, -0.23367080083656, 0.104657779741701, 
    -0.0712098890536212, 0.0300496368530464, -0.118814518160401, 
    -0.0185437691281951, -0.0739127037183073, -0.00187145937111471, 
    -0.216423259707338, -0.00137514998660957, 0.112306251785238, 
    0.265592296107563, 0.203564775631534, 0.0332596394698161, 
    0.242610282543762, 0.544939878561858, 0.348531276002815, 
    0.145897901675301, 0.112276454117244, 0.357147417970655, 
    0.485956715647515, 0.379493840736642, 0.290033833057069, 
    0.302913125229136, 0.327092355012036, 0.281604549274088, 
    0.234976767074986, 0.286878010362498, 0.358437553109084, 
    0.296441813056782, 0.217218310476363, 0.185241971622974, 
    0.257359122814837, 0.270907632556634, 0.157033866253494, 
    0.055430306553195, 0.270920562854796, 0.379995236134806, 
    0.160601858723943, 0.0886702016703757, -0.261064598561591, 
    0.0573095406530276, 0.607557682352116, 0.231504556314203, 
    0.0428067659860541, 0.0028176733768815, -0.307985091572246, 
    0.227136444592488, 0.699789747442542, 0.0647872490786821, 
    -0.028119239442685, -0.262666869798504, 0.363051276788407, 
    0.417294689799373, 0.141483981771059, 0.0214781218477093, 
    -0.15324818291095, -0.141499840550179, 0.430530573426711, 
    0.383550799251378, 0.131831317611733, -0.0480708144482771, 
    -0.0715179831528044, -0.0763887546639814, -0.0743405892106802, 
    0.137604072761323, -0.0946360055216138, -0.011731801907069, 
    -0.140495557630315, 0.134364873386161, 0.10005715210892, 
    0.106136714344118, 0.288894749164569, 0.174210439389969, 
    0.0402417011197467, 0.0252711104745471, 0.239272340122957, 
    0.292398969005003, 0.177525062452163, 0.0746938751060211, 
    0.0122743087998126, 0.166147814104481, 0.218041754903186, 
    0.132875830675747, 0.068462573291322, 0.0421719558064682, 
    0.165118503981686, 0.222712970227875, 0.0953517873466027, 
    -0.00760788646623704, -0.0180038983086778, 0.0395908909903202, 
    0.0194965335419856, 0.0427617621661247, 0.00945118717873551, 
    0.0458331604158575, 0.0136173144974724, 0.0486712394633383, 
    -0.0372235768839636, 0.0941622528362472, 0.108274561553472, 
    -0.00674723762240055, 0.193436542738394, 0.344365435237502, 
    0.123185702348229, -0.00804993508258103, 0.0280363649442325, 
    0.014885926147618, 0.471058207405366, 0.346974080626386, 
    0.0584312010397301, -0.282166699774769, 0.269697022121743, 
    0.553171370114316, 0.198657021625314, 0.0535601589818073, 
    0.0311054027295756, -0.0162736150335758, 0.247540738908229, 
    0.481913826032326, 0.310236357068591, 0.119160290285397, 
    0.129269396544345, 0.106022812919039, -0.0837672525880114, 
    0.113286561020433, 0.0811494422634991, 0.0334715449920806, 
    0.109999747179871, 0.0552950965287754, 0.118513625187091, 
    -0.0534591881923511, 0.108766129251081, -0.0352417804151192, 
    0.106709746465723, -0.246703988657464, 0.0172974457082635, 
    -0.313721255569031, -0.189847646282815, -0.000487955124325687, 
    0.0511603022972821, 0.0761056383931823, 0.0733820685613437, 
    0.0358812282418608, 0.091702576559554, 0.0647966823188237, 
    0.0806609952100095, 0.0248989757001258, -0.0282451823844888,
  0.113995189775337, 0.191017420578575, 0.193400377406876, 0.245964748508451, 
    0.266100492937696, 0.152115920024365, 0.212550673958853, 
    0.504748593639681, 0.277426900175155, 0.0164964986134397, 
    0.0307988562830112, 0.611265461277479, 0.287936096037358, 
    -0.0733593547164391, 0.458571575708972, 0.507122953019382, 
    0.0811833829195427, 0.0381412588511858, -0.270001502669225, 
    0.364232379692455, 0.463216096045259, 0.0652622976561612, 
    -0.140318892899525, -0.123654192447359, 0.499870489271939, 
    0.266304356809604, 0.110611680854347, 0.105791179773384, 
    -0.0663074905418541, 0.669558867212035, 0.131283532431547, 
    -0.0217281460684584, -0.0861429961030816, -0.0479851686277698, 
    0.58098171958069, 0.109339731034092, -0.220494924498158, 
    0.325368888436044, 0.141440558912611, -0.224088148300626, 
    -0.0980401477493511, -0.140981560090352, -0.0961381525176307, 
    -0.147303552370588, -0.141330277313007, -0.174089536251797, 
    -0.0832848418259136, -0.0776535439625529, -0.211820934123153, 
    -0.113582549291496, 0.0190969317110401, -0.138406981133198, 
    0.0714355777520857, -0.107257916548428, -0.00528180213738933, 
    -0.00745401161914147, 0.0682296778523537, -0.103755188472737, 
    0.0638853236710547, -0.145378258374393, -0.0396712453206662, 
    0.0532753110659766, 0.0191000201064332, 0.0327425827479814, 
    0.0364447813189509, 0.0435334680768185, 0.020223578266421, 
    0.0272197690820062, 0.0198739039718597, -0.0496620809430973, 
    0.0441355617345478, 0.183257621612278, 0.147680160408225, 
    0.0364915743351457, 0.097052353048689, 0.333269631265604, 
    0.192631654649294, 0.106237728584155, 0.170430619316704, 
    -0.159331538074964, 0.601897513993929, 0.274171465759334, 
    0.0116223096977184, -0.269613135440135, 0.23420161291666, 
    0.66809748749392, 0.150686742750108, -0.0397440487741435, 
    -0.156511676577483, 0.287982464537786, 0.402666948705027, 
    0.191972721206187, 0.24494236188003, 0.451464158498492, 
    0.0917583962457732, 0.0665695027435504, -0.27229462764198, 
    0.129183163653565, 0.276053225762683, 0.0574008652726788, 
    -0.134133013097618, 0.181162356387429, -0.105326583190466, 
    0.13328419920908, -0.0947155262045345, 0.121706773117111, 
    -0.321985909488778, -0.00299543846342459, -0.290714893198016, 
    -0.208646906638719, -0.0211494915886538, 0.0737525595420809, 
    0.084907117619313, 0.0546559355886258, 0.0771394194986156, 
    0.115181369909827, 0.111962540450071, 0.0729896382629236, 
    0.0510111474945287, -0.00552478325103323, 0.306580699579017, 
    0.198742198711047, -0.0257223732801315, 0.140555017508435, 
    0.398371592965921, 0.3411633355418, 0.18160167865372, -0.138105681054225, 
    0.370580218760769, 0.461245323578794, 0.0843914286548302, 
    -0.15165363585438, -0.116179598384938, 0.616100210118785, 
    0.341356550729336, 0.156381184150993, -0.256977816180271, 
    0.803620544411881, 0.437674394565833, 0.129606994262383, 
    -0.0703470893132967, -0.139581218026238, 0.0642918194964574, 
    -0.119362188171586, -0.0219201341006325, -0.0642810227125472, 
    -0.0166276060825078, -0.0139756077987561, 0.0359612661715152, 
    -0.139181347553321, 0.0187096293697803, 0.222760886667278, 
    0.196690397775784, -0.0131662348922095, -0.0321541004255706, 
    0.580086817538856, 0.4031025072347, 0.115944383111084, 
    -0.054951097073469, 0.110707618418349, 0.387161107224965, 
    0.369861624300124, 0.253415308311224, 0.190759229716311, 
    0.217796776311872, 0.262643012461788, 0.218342821284639, 
    0.167285242008597, 0.225418811874729, 0.277376238102184, 
    0.213134164768911, 0.177785646522751, 0.137429132915467, 
    0.0952499300317052, 0.173663897900381, 0.169150644891627, 
    0.10046953989098, 0.21362417855015, 0.198552390426597, 
    0.0881933627794137, 0.0738748298848052, 0.0976778294656927, 
    -0.286060652743328, 0.429967750078, 0.602767249100098, 0.152045400477992, 
    0.326926967393639, 0.69926171523864, 0.54311676359289, 0.349316279081437, 
    0.200745730420611, 0.135932836779956, 0.136465193445149, 
    0.194856807569606, 0.0707913038784471, -0.0239742026053681, 
    0.0584591836030125, 0.129727851946809, -0.0304183948117638, 
    -0.0377904206480497, -0.0823508896100321, -0.0879765810534655, 
    0.0159878665350734, -0.0736480787895315, 0.0288308771414654, 
    -0.0919849583293343, 0.0156950675685056, -0.0883207421599123, 
    0.00885886428867305, -0.0938956594076123, 0.0233164964582725, 
    0.0126354392597361, 0.206415258297143, 0.154815248929539, 
    -0.00350035776296222, 0.0142349731366124, 0.266616334232652, 
    0.191683572728902, 0.00255847994940334, 0.374564060810609, 
    0.568915836986733, -0.171338398810723, 0.107523928593098, 
    0.818946477409239, 0.278335654610547, 0.164911553985357, 0.2821426222114, 
    -0.09190348256218, 0.256699078587477, 0.896604440775904, 
    0.0744884238110899, -0.0420866631328575, -0.042108428957438, 
    -0.055658621220801, -0.0829056838808388, -0.0938238778610544, 
    -0.0432029055172117, -0.11424694779106, -0.0459088508800339, 
    -0.0928532601672924, 0.0652687806004997, -0.0271954396172724, 
    0.0551800517326392, 0.0183398095077372, 0.0472789107303337, 
    -0.0137158897618834, 0.0429502051620323, -0.0354208319200154, 
    0.00818281133804589, 0.0117112916334413, -0.0119263854765797, 
    0.0709783778121549, 0.174403280914698, 0.115167562529512, 
    0.0521046385140122, 0.0388379287773145, 0.0901645740313169, 
    0.0847022177442979, 0.321501293794863, 0.440137144134388, 
    0.19182675988059, -0.480995865139574, -0.0266870767113632, 
    0.45290872190163, 0.376861445446291, 0.402959797434932, 
    0.0761220866875437, 0.992851724094549, 0.734800877349523, 
    -0.104064131057346, -0.175895051122994, -0.136996476160138, 
    -0.00536551692139216, 0.011405452182714, -0.0782835081348563, 
    -0.0973174415089715, 0.153310466669672, -0.025249289670244, 
    -0.14536972787574, 0.000572996391452245, -0.155038470296179, 
    0.0804144145163884, -0.27079880746684, -0.0624776529094478, 
    -0.0872916642180775, -0.166934639796227, 0.046011144202258, 
    -0.0613268882790079, 0.0779095217509575, -0.192127321632864, 
    -0.0117970188247134, 0.0791884500240529, 0.1141774239023, 
    0.123742636161844, 0.131202284760569, 0.128655946878916, 
    0.114361994291903, 0.115407236531581, 0.16475610812801, 
    0.147291572156981, 0.0945062479128439, 0.0877879626350659, 
    0.0539520046736761, 0.0732900319346004, 0.082607165783948, 
    0.0894154802945038, 0.0593164999644455, 0.0811738065183809, 
    0.0462098248754611, 0.0221171894395201, 0.0699918178529008, 
    0.11227819251645, 0.115106388502752, 0.105001015037046, 
    0.125134907431888, 0.171144254871393, 0.135501017834236, 
    0.0666413378946742, 0.204762957330318, 0.206602979174479, 
    -0.00979871462720179, 0.0414339931007832, 0.403288476344349, 
    0.44989094244886, 0.422929872207456, 0.613194992936815, 
    0.285775204953359, -0.365568060863389, 0.263074731834637, 
    0.386506546049129, -0.0548727983187223, 0.00661717745162752, 
    0.0304433791033002, -0.103169224450337, -0.130244745433438, 
    -0.143072236616007, -0.228617842521183, -0.145375936335642, 
    -0.127087510007171, -0.164596663075785, -0.0695600842105073, 
    -0.174795966582539, 0.0692605599973424, -0.0535824150877146, 
    0.119717359272506, -0.275401299530366, 0.0460967118426142, 
    -0.14759217780992, 0.0154777365082124, -0.323481947545836, 
    -0.0634989724189895, 0.0147540016946161, 0.0468476106727069, 
    0.0764759615482088, 0.0879304942954015, 0.0547869942740027, 
    0.0311859664623545, 0.0800243363077069, 0.0700436542277679, 
    -0.0110269223494038,
  0.113372225720579, -0.110908497134723, 0.0826421899265074, 
    -0.0772734794835369, 0.035036476222725, -0.142758899461405, 
    -0.00495632636527503, -0.0821930800032743, 0.0113047240430038, 
    -0.226496012610209, -0.0352680958242314, 0.0547058878442526, 
    0.0812054443401754, 0.063012642111702, 0.067283243831903, 
    0.0632283826758404, 0.0739723481927495, 0.0790066559722153, 
    0.0683448180229944, 0.0232373255687336, 0.0686682230595673, 
    0.103005915947492, 0.119386475676139, 0.0897433436169041, 
    0.0752779366023615, 0.150240824350695, 0.144537932385009, 
    0.0863419083226839, 0.126085145119324, 0.0648542970374908, 
    -0.184820879768636, -0.0997764697283537, 0.815432709013432, 
    -0.0853547357506706, -0.180698008008877, -0.307477449629568, 
    0.378862658441305, 0.558640634011562, 0.468429563939942, 
    0.212272864091347, -0.234865954872613, 0.119948360399247, 
    0.49589538788541, 0.0894705592336334, -0.0800788601208572, 
    0.194983137879311, 0.252053782783348, -0.057915074505751, 
    0.360997222176113, 0.390760284526364, 0.0595856141386224, 
    0.0249879817007444, 0.0236912799995947, 0.0221548238664588, 
    0.0244422316759127, 0.0237893859346347, 0.0226751352798517, 
    0.0490422317639134, -0.0359947159975744, -0.00121818539266853, 
    0.446442938880067, 0.0780373933447339, -0.108414427074832, 
    0.0619143944849479, 0.479367913591691, 0.422401096901136, 
    0.266148805432691, 0.142547345699, 0.0151848505307396, 0.756002555629189, 
    0.375938364738237, 0.108205025807574, 0.225347864190227, 
    0.372989486326104, 0.147393894685449, 0.796649892532593, 
    0.580295128356189, 0.210059850966623, -0.0461342698935125, 
    0.544249543910293, 0.353043561689904, 0.147848759047928, 
    0.135238062888113, 0.243225159492667, 0.0982771042031382, 
    -0.122744444276851, 0.0150411381106075, 0.257121066876676, 
    0.27078702908268, 0.130658414463713, -0.169193690376126, 
    0.13329662063498, 0.340420045571988, 0.0256570015744268, 
    0.407977940976419, 0.339782610378218, -0.000822102667959373, 
    0.0202946565921217, 0.0966924438741145, 0.0279946390100417, 
    0.0602307194751985, 0.473987960848496, 0.182266416733441, 
    0.00436613479699535, 0.115999051730673, 0.25834924523522, 
    0.0665155747705878, 0.21396489960773, 0.391239798706074, 
    0.0106712272411079, -0.0992517800113796, -0.0032233124551999, 
    -0.105275948886614, -0.022825724578404, -0.044205267110826, 
    0.0106115427528093, -0.231308848432064, -0.0208327483451789, 
    -0.181380674742658, -0.197485280939703, -0.0217331697537675, 
    0.0933093588172235, 0.284405578459669, 0.173972096846505, 
    -0.0259653523181588, 0.0126199836909939, 0.452382493874287, 
    0.335880191458824, 0.139725622410497, 0.0668530621623907, 
    0.177953123916678, 0.197590122680529, 0.222848037365362, 
    0.486582471215779, 0.532076800561218, 0.335709703281431, 
    0.274414901785055, 0.385236535599527, 0.302861378473698, 
    0.23110829718212, 0.486048825294693, 0.47265628476019, 0.231478264812062, 
    0.139657961117605, 0.149045775319772, 0.193752039652923, 
    0.568181950419617, 0.440685626620552, 0.081745278059558, 
    -0.133730546137425, 0.0426359837370567, 0.236196181253464, 
    0.629069485107059, 0.473210932272548, 0.1120569474807, 0.13041910314353, 
    -0.147657239944727, 0.862819891721274, 0.105794053427544, 
    0.014237261531519, -0.169503335912636, -0.180194848875227, 
    -0.0541833795665639, -0.214112051291485, -0.0943879976111289, 
    -0.154772897626701, -0.0848248164351199, -0.158828545233339, 
    0.0195346542922171, -0.166567255585564, 0.0670328351666458, 
    0.0531197644595627, 0.0729447693131255, 0.0734192735055442, 
    0.0811536229272033, 0.0492052532215749, 0.0726341660649569, 
    0.0594693133033351, 0.0684364753497561, 0.018083292006203, 
    0.0526834504967215, 0.106315232021562, 0.114953244157551, 
    0.161462541383659, 0.128256097933185, 0.100686915795718, 
    0.309274650743482, 0.155644901677382, -0.102048745070013, 
    0.0200476760136184, 0.488470796810371, 0.224557704052285, 
    0.141499578747071, 0.111251048655687, 0.85631997836411, 
    0.150707182614878, 0.0855865745901686, 0.553651213926794, 
    0.0775307358169505, -0.0134366687690459, -0.109183956342565, 
    -0.180746983403174, 0.00235053672145817, -0.184123449192898, 
    0.0724954563796696, -0.167180528338707, 0.0786542232121655, 
    -0.183608825863767, 0.0379240641852439, -0.0659798920956251, 
    0.180692277504167, 0.00915674174672558, 0.0701334026255365, 
    0.0523887319258334, 0.087823561212941, 0.046830498758016, 
    0.0835091169101535, 0.0352753437804225, 0.0530018986166361, 
    -0.0703439310904388, -0.00764798384341389, 0.0225231909881754, 
    0.0181615875870477, 0.0227837808340309, 0.0346460070231931, 
    0.0144872253942421, 0.00967710082694571, 0.128438211222979, 
    0.0857610867273208, 0.0213596414710413, 0.542376837431741, 
    0.0673102736146704, 0.499899811468579, 0.655147911038076, 
    0.173328245236077, 0.0354701831106697, -0.122747967004224, 
    -0.148532197140656, 0.676206896214788, 0.511204189083572, 
    0.245310527389824, 0.238773678165089, -0.237305696033262, 
    0.435879117724398, 0.225989491555315, 0.0242781330835744, 
    0.14404640645464, 0.411145547381893, 0.120035419366583, 
    0.186985085586675, -0.231959880287469, 0.234737717793405, 
    -0.151084766138463, 0.122883224402636, -0.454015419931687, 
    -0.0719635508289889, -0.113915556194785, -0.165896240626613, 
    0.179259893882796, -0.364368979297979, -0.0445853330857615, 
    0.0896064083162014, 0.147612015271234, 0.151559172763809, 
    0.155673669601781, 0.122923467955107, 0.123367351962829, 
    0.12227607762412, 0.144024688267324, 0.158990022520153, 
    0.0972748061034051, 0.0762283638269384, 0.0260855742020341, 
    0.062746534232386, 0.0380335126955702, 0.0205202840743547, 
    0.0428771306529015, 0.0922064510982685, 0.0934635599856531, 
    0.016480038242916, 0.0810206491936532, 0.136694981600233, 
    0.105620262745232, 0.0619498994844455, 0.144227440110462, 
    0.294757123438999, 0.134674157933831, -0.00779499846785124, 
    -0.0722570197990787, 0.0606122471884681, 0.500898793199598, 
    0.282956848165154, 0.222020875079844, -0.312391484837087, 
    0.621576386881553, 0.415051211809958, 0.18893896355901, 
    0.0583548590163212, -0.247836272660042, 0.00847838866304072, 
    0.377684503550736, 0.258616847878131, 0.480750877161967, 0.3670931577905, 
    -0.0506147484653753, 0.17796554789927, 0.206049797562519, 
    0.449801446543726, 0.291492926163838, -0.126029916830798, 
    -0.239389124848888, -0.0408599379027257, -0.334621631783573, 
    -0.210141258713843, 0.0525984876670435, -0.219050650929312, 
    0.0630374372182998, -0.153246499795755, 0.0262904722608305, 
    -0.260337667334906, -0.0180240452068564, -0.0201007772042523, 
    0.179795562964382, 0.284105530673181, 0.142257412739257, 
    0.0672155891285597, 0.0608685959788934, 0.573808465211158, 
    -0.204764369246617, -0.205834439848274, -0.116061184301074, 
    0.734490931574701, -0.0124745746727981, 0.0263567213161006, 
    -0.354221918459716, 0.735388182953912, 0.418240530703665, 
    0.170613375081569, -0.257435325973392, 0.303407367872564, 
    0.511019385616343, 0.102777785790306, -0.142950718669402, 
    0.047480791058196, 0.217050374273793, 0.359230555907627, 
    0.25318046327742, 0.0575412636339718, 0.408687544273932, 
    -0.00859658013427601, -0.152269347833953, -0.21976852181097, 
    0.0372891220604133, -0.176482193585147, -0.136518098966369, 
    -0.206619780205679, -0.0393692615928858, -0.315082445915506, 
    0.0561454622500438, -0.159027325340036,
  0.0644190618231183, 0.0770969480645376, 0.0548489844611934, 
    0.0656362102119261, 0.0559907876768974, 0.0573167438669733, 
    0.0448737593226016, 0.0839689111380271, 0.0454248797870436, 
    0.00459354010909623, 0.322249017354105, 0.185235064006033, 
    0.0622091492202482, -0.0866399535357645, 0.490775321329575, 
    0.216305843692862, -0.0266580587520728, -0.181135020591558, 
    0.300120092805031, 0.470804078905622, 0.593542125059426, 
    0.298094536042882, 0.0795156870387749, 0.0561370764546239, 
    -0.240666148295046, -0.67683214462142, 0.414919581466858, 
    0.625318987893339, -0.118811093445193, -0.228799346290016, 
    -0.154923195351077, -0.29247127536598, 0.0233867015257469, 
    -0.341987026420052, -0.135417546699319, -0.27703747088777, 
    -0.2608310343685, -0.141960780569187, -0.270245285516045, 
    -0.136785207001833, 0.00641021575588487, 0.122161383391892, 
    0.0982479449484179, 0.138201465123106, 0.0349373749966491, 
    0.0906119316906967, 0.0652958034959174, 0.0923431945453232, 
    0.159429143831746, 0.0753001225666765, 0.0735474876092166, 
    0.0694688583186823, 0.0783710081246717, 0.0762962464638083, 
    0.0926167211018368, 0.0708924318857006, 0.0861905399240794, 
    0.0726307905941327, 0.0863977577549289, 0.0397828530526644, 
    0.0872509506023425, 0.113183854033283, 0.114501021260394, 
    0.12309356510091, 0.150231102044956, 0.121681275225933, 
    0.0585784692374488, 0.119420055536999, 0.201827222602892, 
    0.170674339116505, 0.182043789668198, -0.107753675705388, 
    0.43784318227546, 0.306302718637555, 0.068982826735852, 
    0.00280340463459888, -0.0336776587547019, 0.743093189674401, 
    0.164684802789262, -0.0948376259645674, -0.208587660170981, 
    0.321871184099741, 0.680572080484627, 0.0382605894296154, 
    -0.193462864609329, -0.195571024010938, 0.477135516509868, 
    0.269735342642545, 0.212598232342147, 0.267530134654525, 
    -0.136563809083145, -0.268633170813574, -0.116220491723924, 
    -0.197381061067502, -0.123662886656294, -0.20473241401815, 
    -0.142235545474204, -0.173318735655806, -0.0400966292188335, 
    -0.30626984462121, 0.0673466420762994, -0.136286411477322, 
    -0.0523530215434281, -0.0863266836532238, -0.0748403547854127, 
    0.0131603665112135, -0.0717461049346932, 0.0939983222128366, 
    -0.0740152065318638, 0.0556432160159663, -0.0201470599502099, 
    0.0404448004552442, -0.0353693002885324, 0.0107760594757583, 
    -0.104599386886466, -0.0247166779638229, -0.0150461863792444, 
    -0.0129165211197176, -0.00296800112224904, -0.0845746941262338, 
    -0.00986615052862769, 0.0682494417892975, 0.078356162038149, 
    0.0304362458951719, 0.0475630341890629, 0.175381543540029, 
    0.0859878480182594, 0.0858758504524118, 0.25474582806789, 
    -0.210316214292444, 0.498600859259045, 0.336369600809269, 
    -0.00805922579208911, -0.119182234484752, -0.0707288253177219, 
    0.595008097366794, 0.364125853009, 0.322117705404808, 0.758781986250404, 
    0.388256094733139, 0.159388520756043, -0.435838561744154, 
    0.369053911136604, 0.330535081209942, -0.0368152273330052, 
    -0.0394646668017701, -0.25217349231337, 0.517490343212178, 
    0.210475815809202, 0.066773909253852, -0.23225137746961, 
    0.084076268535263, -0.319067693016369, -0.100588884186951, 
    -0.213495430766231, -0.211557959750283, -0.0506277105838775, 
    -0.214669767131251, 0.0655942325718823, -0.250003094032744, 
    0.0436232185353737, 0.11838835768037, 0.092782383109663, 
    0.0845961227451533, 0.0716503572005113, 0.0841703477209916, 
    0.0967366855532103, 0.0858383446888956, 0.106846894212357, 
    0.107960875400323, 0.0443660406093324, 0.0550203360040803, 
    0.0557295853635004, 0.0610678614089056, 0.0394472764262492, 
    0.0628940789414821, 0.0358410051272246, 0.0480443878669397, 
    0.0259528906442355, 0.00389801653911274, 0.0559411240917003, 
    0.101271933011078, 0.111330672066821, 0.124891511631255, 
    0.135216240064846, 0.0963710378993136, 0.0799977504616373, 
    0.189260132665466, 0.149584123505676, 0.0730130801612908, 
    0.0904934551946417, -0.063787214305998, 0.383755594559522, 
    0.355254172042824, 0.00634589983081937, 0.122755721224542, 
    0.70936398921078, 0.238451379596544, 0.169095876178419, 
    -0.0642805267138424, 0.605475490725903, 0.183161357819459, 
    -0.00540582415814461, 0.428848392094471, 0.187912777762324, 
    -0.0866206639344812, 0.0263150258499683, 0.204703086724355, 
    0.675674840001247, -0.372098621128524, -0.119366591255787, 
    -0.296973063140725, 0.0393148124155918, -0.293855915919907, 
    0.0228128819730224, -0.375759551914912, -0.0715201078478503, 
    -0.261059424920608, -0.0826918009543949, -0.25687260664711, 
    -0.0109750125111801, 0.127089761688146, 0.0542022892370511, 
    0.0680727196412741, 0.0134748319077549, -0.0434695521041807, 
    0.0986143332816362, 0.104205726944402, 0.110639512754873, 
    0.00812851254380054, 0.0312925098489435, 0.0718413597657751, 
    0.0768136804616444, 0.0712064741558153, 0.108520586443104, 
    0.0988969154167565, 0.0467230676642928, 0.110856326740853, 
    0.241736165825265, 0.151951615775576, -0.0198467095790461, 
    -0.0479210943107057, 0.626610919543748, 0.237102170958356, 
    0.151968012695255, -0.300343148768746, 0.368057932520483, 
    0.419728187971538, -0.150367643602354, 0.323946600665216, 
    0.890829630444062, -0.0941879797824041, -0.290321065550444, 
    0.419540172272201, 0.304422143223975, 0.0896752347372809, 
    -0.254527194516077, 0.26817143328116, 0.122589673519622, 
    -0.1688287628542, -0.248338889232464, -0.190728282424796, 
    -0.171430317367133, -0.224165687294344, -0.0804121706841542, 
    -0.230496041953647, -0.0949694745310265, -0.128492821705194, 
    -0.12473839583825, -0.00843049811995098, -0.236113540710862, 
    0.180216304311434, 0.222978661411026, 0.078443246228888, 
    0.0605342040394571, 0.118674521085152, 0.322414267464357, 
    0.207210327959291, -0.0804397087275576, 0.355658255156813, 
    0.682065862938017, 0.431692873704795, 0.264299027745085, 
    -0.294031591096212, 0.957165032384933, 0.718472667185008, 
    0.259804216601649, 0.120253946766602, 0.9157859416494, 0.226221200238138, 
    -0.0927113995446799, 0.0401121761156185, 0.0367345695819581, 
    -0.272172534028053, -0.021023409990306, -0.124920348816938, 
    -0.133068615850804, 0.0741723011475735, 0.020817135269694, 
    -0.186478355011322, -0.0616285039396401, -0.0632189334962016, 
    0.0465685463040528, -0.162764800260657, 0.0117391492501285, 
    -0.142069858612855, -0.0827687071963627, -0.0725577657060669, 
    -0.0302020090307244, -0.0892545735234873, 0.0527447767401478, 
    0.06515956733183, 0.0881386837470405, 0.110507991982961, 
    0.105507131712193, 0.095404640285716, 0.0788278895672649, 
    0.0776495102179151, 0.114727850873928, 0.115462985572852, 
    0.0575588656879418, 0.0276438980922026, 0.0464304059348804, 
    0.0487800988681413, 0.0580252724238184, 0.0221744646420509, 
    0.0448149953674098, 0.0625658060742014, 0.0717056247001182, 
    0.00695631278220254, 0.0720093999364348, 0.0800601374514642, 
    0.109083413946126, 0.162109074087295, 0.116576423630351, 
    0.0104561299963442, 0.284697823101825, 0.174699036420327, 
    -0.142875604124122, 0.0452426131283091, 0.586187110553762, 
    0.100018879700252, -0.167322039225715, 0.558948121574708, 
    0.367522411008543, 0.24496618565049, 0.411486171961172, 
    0.212460968112618, 0.395722060614547, 0.874212989863371, 
    0.151094412885101, 0.0177990590775155, 0.0156046213318323, 
    0.0146602088928128, 0.0267450451091572, 0.0114138065929828, 
    0.0415607500053483, 0.0229545229964759, 0.0219092552777099, 
    0.020042488450746,
  -0.200625582848237, -0.0544356562471925, -0.25055880354169, 
    -0.103357903310361, -0.195278383702156, -0.153711710140969, 
    -0.153518497664521, -0.16856951501688, -0.0559239010843818, 
    -0.194839342733148, 0.0307256802581942, -0.110403105915601, 
    -0.0316993834994347, -0.0332189905849001, 0.0106169577143135, 
    0.0170163321403107, 0.118229912880557, -0.146175946793306, 
    0.0936678032617948, -0.0685757939686637, 0.105656472082213, 
    0.0186538859102306, 0.129768580417009, 0.160813470923962, 
    0.100889752098401, 0.174445791724552, 0.121323288574356, 
    -0.0102726552468329, -0.301807045034163, 0.484091753755597, 
    0.384494167145973, -0.224193518478599, 0.205352298884471, 
    0.60876514238757, 0.00724066318032808, -0.0904275269759352, 
    -0.249604970901784, 0.650857020839751, 1.03102999216285, 
    0.122785545544577, -0.211967480057113, -0.0958739241307254, 
    0.231749252245314, 0.269206431296534, 0.155577276475104, 
    0.00587482555179852, 0.413010967263261, 0.0565629603407824, 
    -0.172353909262759, -0.105866429392859, -0.103352480678782, 
    -0.255395279535584, -0.0170784191782408, -0.24853777127507, 
    -0.0565505296827323, -0.215078703678554, -0.0478839438954327, 
    -0.18249885483593, 0.0195115316072321, -0.205417702785062, 
    -0.00916772320940405, 0.0489358811123724, 0.0619514034925319, 
    0.0648113862320498, 0.0636702618004265, 0.0620110974695619, 
    0.0691616338970112, 0.0840321770176767, 0.0693821914620199, 
    -0.146148632893183, 0.217671906625225, 0.405287029954854, 
    0.205875995093107, 0.168674526568715, 0.873993605518101, 
    0.258924676258337, 0.080504075457905, -0.1957517379632, 
    0.151298508607204, 0.721555254111704, 0.112133374916629, 
    0.0789576516744605, -0.463194145684974, 0.0430621546755479, 
    0.629446889913119, 0.237814439207047, 0.0432703082718772, 
    0.0981765597197945, -0.167848899375142, 0.365959336068785, 
    0.583424271317204, 0.202877403939449, 0.021010550130985, 
    0.0212923627377156, -0.0447622933367161, 0.118462679212739, 
    -0.0164479592811065, -0.0407907168038798, -0.0886587537961971, 
    -0.0546802173918088, -0.00663863880553745, 0.233746538594382, 
    0.381954846149839, 0.132198171973591, 0.00930641581545265, 
    -0.0866130160624089, -0.037068640503625, 0.318427265917185, 
    0.333046057804146, 0.123275919412092, -0.000294620725829017, 
    -0.0483802779516649, 0.178614660924409, 0.102317307133487, 
    0.0510609877098251, 0.0406899580436893, 0.0759696496578035, 
    0.193025673069568, 0.0992348360582003, 0.0382568159934875, 
    -0.138176947990187, 0.0429060390759078, -0.16003931370635, 
    -0.0739820960455308, 0.000461662320239129, 0.0850913573250662, 
    -0.1011634160382, 0.10615380931609, -0.28368713668472, 
    -0.0775383520866834, -0.0426042591884118, 0.0446199293996157, 
    0.00815582394287162, 0.0470799754716445, 0.108188279436789, 
    0.0931494097090474, 0.0708335214735868, -0.121948149965786, 
    0.0348556574909465, 0.266619859089343, 0.113399621057407, 
    -0.0901318767215337, 0.0231932073174532, -0.0287447453023354, 
    0.913725110557247, -0.271876021404397, -0.650470878441761, 
    0.266039331134371, 0.438520294015012, -0.308686355169135, 
    -0.123060810657654, -0.113694587792032, -0.0104808510344327, 
    -0.159582976908596, -0.0278775117453357, -0.069796777618647, 
    0.041387809794807, -0.0999323917333301, -0.0805341470467365, 
    -0.082872452773403, -0.00821337552503868, -0.150263061676763, 
    0.0199272043120362, -0.0773151436927579, 0.0168031810973825, 
    -0.168362359491825, 0.00203738336906911, -0.0642493584421452, 
    0.0395689421711121, -0.213846580731041, -0.00938707361421871, 
    0.0559713303205453, 0.0646338709470379, 0.0740351935160262, 
    0.0777617545353482, 0.0590144127133867, 0.0698869432913297, 
    0.111234863451914, 0.0737738602903645, -0.00114793728959171, 
    0.150285640366544, 0.184486481807915, 0.0906196629381943, 
    0.214792950108898, 0.352524546022168, 0.168732731186003, 
    0.00760709845786337, 0.324396669533908, 0.458204227375153, 
    0.199266162528209, -0.134406722607869, 0.44980924810713, 
    0.331760496222187, -0.0494230303078035, 0.0968642093030294, 
    0.642379285858958, 0.229507321005121, -0.127105497947957, 
    0.528588476091519, 0.402199539576961, 0.0363920318837219, 
    0.0357187517233052, -0.100389352926171, 0.0805472041647118, 
    0.0471088609536411, 0.0934935356865912, 0.179271947676509, 
    0.679881426208794, 0.12774903683829, -0.2157422135552, 
    -0.272409897743549, 0.0109163777232969, -0.241658008315625, 
    -0.0893336420695894, -0.195977249770487, -0.151017785338928, 
    -0.101188324455863, -0.160885114720771, 0.0202538877901554, 
    -0.167697445537059, 0.0970769865697594, -0.00278700902981471, 
    0.0512931121390644, 0.021032685986038, 0.0531808926107443, 
    0.00717031718489994, 0.0497998475274168, 0.037745463805223, 
    0.0523423087880429, -0.0443422889171069, 0.0320948572946904, 
    0.115091851661572, 0.0568964359966817, 0.0797278384052489, 
    0.149068152281416, 0.231034717537059, 0.170180572883649, 
    -0.0541908311596017, 0.26717537790552, 0.166982795001067, 
    0.191228687857769, 0.321366207183979, -0.123963292357962, 
    0.919672815909933, 0.357350461009064, 0.0595723343383058, 
    0.081177782501537, 0.180131462460244, 0.0145756265470133, 
    0.712355315095949, 0.522010727240049, 0.1199768461763, 
    -0.0397349222832692, -0.277411613740463, -0.00512962907453216, 
    0.0702704574229151, -0.115270924135076, -0.0339015974395638, 
    -0.0689469580011433, 0.0761658397155143, -0.361409186033841, 
    -0.0657177948824171, 0.0142815082722738, -0.198035238436319, 
    0.293209796558993, -0.233237767321411, -0.030834620199134, 
    0.00193937145310687, 0.0802085457935689, -0.228008085792036, 
    0.0543235868771441, 0.0367769255278989, 0.0396281160854747, 
    0.0538072627348691, 0.0597874988448239, 0.0437599220449391, 
    0.0561326338804783, 0.0607750882509596, 0.0490088250237283, 
    -0.00565535587879161, 0.0600252369249765, 0.0955620534921679, 
    0.16745875774141, 0.137140669293666, 0.0619273616703153, 
    0.206789841944189, 0.248240486632361, 0.076469557201574, 
    0.0412011569117072, 0.239897758285684, -0.0159508688574173, 
    0.752518045729083, 0.237469836832077, 0.090514157030749, 
    -0.391715438035839, 0.244927197760941, 0.692971158106176, 
    0.258108652209927, -0.107913174507393, 0.307419326113487, 
    0.213289456071334, -0.0500308121379717, -0.110077026741962, 
    0.0512371629991216, -0.00566152133345083, 0.00282546671610838, 
    0.00517520711708799, -0.13109430823812, -0.0377087997323909, 
    -0.0960446279605167, 0.0361114705160366, -0.308381961910028, 
    0.00598553738852821, -0.0918641497473315, 0.0289370604382207, 
    -0.184001028987766, 0.0420701845505344, -0.0912121326116735, 
    0.064302036809198, -0.301606951096445, -0.0110433669186003, 
    0.0561043137934675, 0.0578580260470462, 0.138389395131419, 
    0.185715660975201, 0.116061378032705, 0.0966959888848715, 
    0.254146078054239, 0.192215015189619, 0.0240993635807734, 
    0.363945068843716, 0.449916642479993, 0.171884316723912, 
    -0.0783436581118951, 0.711400122001689, 0.334337631216192, 
    -0.0203740440734266, -0.0439313592978561, 0.734301109145985, 
    0.301872273304243, 0.0676320993806278, -0.0168896316973101, 
    0.0980700437592737, 0.0322178777337477, 0.634999998532313, 
    0.580282836837445, 0.0359254183647646, -0.0159000071434504, 
    -0.260511046120943, 0.403499161209761, 0.298758991837563, 
    0.196372958651049, 0.188712037458948, 0.374640269045386, 0.3014643949583, 
    -0.149588852287606, -0.30724483303221, 0.188848867394678, 
    0.0056129587979584, -0.21115755458323,
  -0.052589935153911, -0.241414366872108, 0.134958079029185, 
    -0.0634865168000007, 0.157516726178341, -0.0925590611428011, 
    0.160131843232209, -0.203246037559717, 0.0941092731419159, 
    -0.289878744350803, -0.0313633603482177, 0.0406868468490461, 
    0.102837045807583, 0.139217134934157, 0.0958861642490277, 
    0.123002821949582, 0.252269019919239, 0.0946231026296729, 
    0.0269581290436817, -0.106147013337843, 0.51931969890802, 
    0.0198082938467312, 0.540627795859868, 0.720072688945183, 
    0.0435078329699065, 0.0810005001506226, -0.0941383056691016, 
    0.0101543979023722, -0.0155413612762882, 0.664883261219775, 
    0.515768717673576, 0.132582466494506, 0.0137296760347958, 
    0.0345828819053414, 0.0950878597383826, 0.00440400764930288, 
    0.0599126203358867, 0.125580006825386, -0.0379765158525312, 
    -0.048420323467488, -0.0156553555615884, -0.11756949436189, 
    0.034002283822126, -0.0472584453610814, 0.0462302942437402, 
    -0.111458634104744, 0.0416471193678129, -0.0876863386358795, 
    0.0184669067633938, -0.144267504964776, -0.0214030712418555, 
    0.0158972810594169, 0.043610522147977, 0.0377393092575665, 
    0.0143284184396803, 0.0130140989992783, 0.079299750665465, 
    0.111216148305112, -0.0524632037095554, 0.0487046701100734, 
    0.637975898585616, 0.0457466583123231, 0.372605839136507, 
    0.389037088615004, 0.321393917003028, 0.79730474811678, 
    0.338768098448717, 0.0293225984012407, 0.139221671131515, 
    -0.16614502661865, -0.191318781121754, 0.236083308886177, 
    0.343207950908488, 0.354646199806906, 0.470788298789307, 
    0.38373715199464, 0.198813983824922, 0.230998549061495, 
    0.484416404800171, 0.33034710439519, 0.0974951782395123, 0.3260798514394, 
    0.417770937395109, 0.0688260614998237, -0.0825741963427317, 
    -0.0284112863957863, 0.312029048719112, 0.280604207059861, 
    0.254841032190886, -0.138792342267272, 0.489128998395324, 
    0.280129915199677, 0.20491608022377, 0.266643723211762, 
    0.0539632179519542, 0.759648958570804, 0.142719589705618, 
    0.0123778103363186, -0.182969507777803, 0.499855814039651, 
    0.305717140486395, 0.151307454199292, 0.0994399783504637, 
    0.119914876133453, 0.200887371854541, 0.0195645791660152, 
    0.345570614615507, 0.286411000766583, -0.0585858136000524, 
    -0.0666804748270677, -0.336101112322084, -0.112562045779183, 
    -0.111911004673007, -0.223409644289236, 0.0695448323638857, 
    -0.211614544437477, 0.0795573113860139, -0.174665365943892, 
    0.0633513373691733, -0.21806104195104, -0.0107847561456985, 
    0.0657668457212316, 0.0912791435068955, 0.164616017019198, 
    0.20348074835629, 0.131471743242553, 0.114428900212867, 
    0.266817328395172, 0.218238557697099, 0.145422464329597, 
    0.185864137490052, -0.159430812558185, 0.28464649710167, 
    0.677680408644229, 0.0929657437771085, -0.00526158196019312, 
    -0.274627783861869, 0.634781444801134, 0.340321844914073, 
    0.0244306618215394, 0.580158406620455, 0.486072905662563, 
    0.211946590789562, 0.098416509060818, 0.369808737328592, 
    0.502001471818277, -0.335396231733513, -0.0402739855029576, 
    1.01431743697507, 0.195634916033619, -0.0219639092044242, 
    -0.00450778699273634, 0.185161047113949, 2.43903951400448e-05, 
    0.24843021142424, 0.0926305271767095, -0.0672809678349976, 
    0.0791291673958598, 0.280531181162351, -0.0493184078014048, 
    -0.032829350049964, -0.0381460450891291, 0.0139592551703851, 
    -0.0373653197195567, 0.00671082500256598, -0.0520113275478915, 
    -0.0387794280587853, 0.0306566328081304, 0.0354872078769226, 
    -0.0466580217782817, 0.23853923719714, -0.148334236170519, 
    0.206805314597396, 0.372208121187578, 0.333209775839451, 
    0.27778743854837, 0.0310825900435679, 0.719455738659269, 
    0.0380595493162972, -0.0544167110945992, -0.443408034113441, 
    -0.0303551386738356, 0.898506406129937, 0.0571965398878861, 
    -0.0396120920423673, -0.345916029939977, 0.468228460846129, 
    0.54826063225931, 0.290467701903689, 0.197859858757515, 0.16068473927259, 
    0.227849231436137, -0.00307321291534932, -0.0467074332472719, 
    -0.142079517454797, 0.0302898184673765, -0.116191974255534, 
    -0.16354401659302, 0.0122635438262817, -0.14819078931864, 
    0.107090513660638, 0.0707296201050393, 0.067999143900539, 
    0.0450763516573713, 0.105217890930082, 0.0755409158047059, 
    0.0419483066466005, 0.0773515365301212, 0.0913451321836, 
    -0.0187351514222385, 0.149879552277644, 0.23725797575572, 
    0.118959268013505, 0.148570491354064, 0.365462342379946, 
    0.206168714073538, -0.0135353497584881, 0.269260540689932, 
    0.445876257116394, 0.04721050617984, -0.249434414455178, 
    0.0386114022817289, 0.641832985866583, 0.0699645673697976, 
    0.00378648771386109, 0.0912800370000022, 0.0843783465373561, 
    -0.0761789985757011, 0.541822005757333, 0.468555006546461, 
    0.264426601739969, 0.528455937199398, 0.350590333489546, 
    0.10165237164872, 0.115145755378295, 0.309637845853093, 
    0.0982840700662783, 0.0224982560932146, 0.442996842354969, 
    0.19469462838116, 0.0254817157226836, 0.0183087101923487, 
    0.0410201616017602, 0.0430074738236163, 0.0566676892848233, 
    0.0468030614928822, -0.0468248822608633, 0.164704861333033, 
    0.110800570809472, -0.152117102458252, -0.0187700496355886, 
    0.371592323498148, 0.259173037004076, 0.214258142448688, 
    -0.238139442743955, 0.372075909601275, 0.459685274978763, 
    0.150978119467839, -0.20192358314422, 0.138040369793372, 
    0.441807833791676, 0.187288188829179, -0.00203167835690597, 
    0.430705361093147, 0.299246796950777, -0.0933421127260129, 
    -0.306399196372508, -0.278482003620395, 0.628505682695339, 
    0.0680429687702565, -0.162956065093351, 0.163252819804177, 
    -0.0719790031459039, 0.0482508575717315, -0.0811672070064921, 
    0.113451448228741, -0.330326704079448, 0.0237095434215769, 
    -0.372680010108548, -0.209945193955816, -0.0350594446843956, 
    0.0877494573054324, 0.183375397531314, 0.163001321059595, 
    0.110281853677779, 0.11980260327267, 0.0735827416700572, 0.1500481701604, 
    0.21808933902743, 0.153819835672148, 0.125678985095219, 
    0.127801722314968, 0.143665106459168, 0.168894427460584, 
    0.173715274023438, 0.146382304777952, 0.133272066578897, 
    0.160194457394597, 0.160508576650214, 0.134353355209804, 
    0.14596375453409, 0.158615554506355, 0.177145157133625, 
    0.213970158566472, 0.209107480053685, 0.120438556729944, 
    0.0481174047525794, 0.503384407223185, 0.250007889765861, 
    -0.375148534434695, 0.262260823712598, 0.57102814927578, 
    0.0708889905511087, 0.0289618217007124, -0.0991039909777302, 
    -0.438075531398474, 0.487465997968808, 0.374600294061071, 
    0.261674957278068, 0.625706178116032, 0.113694495354964, 
    -0.152405204093098, -0.0949662312759174, 0.625873205241986, 
    0.15428478822803, 0.0876130910416168, -0.124702638428854, 
    0.0253294246117965, 0.311037802176647, 0.324292886137273, 
    0.209960676962456, 0.142436543836619, 0.0575755442947438, 
    0.167431645587864, 0.257205288788205, 0.127162430160284, 
    0.0267681095985185, 0.255956901988382, 0.261317483009013, 
    -0.299625214862556, 0.273593721395124, 0.348306315650476, 
    -0.00872511147853529, 0.377718606077837, 0.436841041603787, 
    -0.00922220960601944, -0.122798796976749, -0.0916524379423273, 
    0.626729540256039, 0.0687546097424706, -0.0390629937727344, 
    -0.0215384796118618, -0.160940110987194, 0.341003593101185, 
    0.228169392248204, 0.397125530284499, 0.591225262450785, 
    0.112698244248612, 0.00647258452981661, 0.0761116143582774,
  -0.17011588848661, 0.320586022384566, 0.2615058009415, 0.22220499158542, 
    0.800948387698097, 0.338113361313597, -0.00843139869244514, 
    0.349082926287057, 0.457967086203903, 0.291680578654049, 
    0.290396708664343, -0.270044456348131, 0.175995178744188, 
    0.480968569897983, 0.29620166271116, 0.0633718795138168, 
    -0.0220441241712361, 1.13782480987716, 0.121945881737219, 
    -0.0543220589116172, -0.156079890493104, -0.10470204094343, 
    -0.132923878234649, -0.128818020653485, -0.0955903631267153, 
    -0.135678180124018, -0.0488977122780568, -0.12887768888729, 
    0.0147385382358243, -0.16639701441341, 0.00463350627341097, 
    0.146921103373945, 0.155138407021558, 0.0961798818569233, 
    0.0881242019726839, 0.310344829437024, 0.391819037762216, 
    0.158795244928963, 0.03082769504186, -0.144864172785029, 
    0.731137906920763, 0.163514176102844, -0.16814569726025, 
    -0.00441904596899694, 0.612927664109725, 0.406889614274836, 
    0.245132979463206, -0.253187876006393, 0.439294702909085, 
    0.451562949799258, 0.303650728192853, 0.194369443902622, 
    -0.164716822991405, -0.0410835192946967, 0.719345210522274, 
    0.146182255815834, 0.0746597762226399, 0.132984905944864, 
    -0.26232812933989, 0.199789065099897, 0.437006481085462, 
    -0.0530321972124039, -0.109252684894532, -0.0500783440300627, 
    -0.106696615277025, -0.108485463494002, -0.146222027734168, 
    0.0357898638201405, 0.201015236679839, -0.133938620935836, 
    -0.171765114102144, 0.0137020992215737, -0.178896617640984, 
    0.00385502898853191, -0.21255789577113, -0.043468369882945, 
    -0.149770267425937, -0.0252334691878896, -0.131208342441276, 
    0.0139137196857073, -0.0632504229869112, 0.0401296806026807, 
    -0.101720340635277, -0.0231096058119508, -0.0229095412202408, 
    0.00195500597075918, -0.101586192070099, -0.0457184989294643, 
    -0.0973868709045745, -0.125442986255658, 0.0257657426114471, 
    0.125606638709856, 0.00753144295460038, 0.0861810683052717, 
    0.252798907369261, 0.0421263671006301, -0.0599628715617558, 
    0.0976292469720938, 0.2490370603556, 0.000533415258670081, 
    0.323871936125423, 0.251914775528978, -0.0808838087982783, 
    -0.395571726412179, 0.208022070740212, 1.16192494757719, 
    0.28458294971408, -0.522738158023502, 0.512596322740352, 
    0.580745706084152, -0.0387491145792823, -0.0799590228048247, 
    0.181328894093987, 0.107132098325374, 0.00650690133681467, 
    0.0922045562195367, 0.110121087533468, -0.138056824578143, 
    -0.163236815218936, 0.0886755408645488, -0.341124452120437, 
    -0.115042686523291, -0.11934047330571, -0.211605546718939, 
    0.0482610477140732, -0.16095651444728, 0.105052243328412, 
    -0.118444351713978, 0.118753949447779, -0.196669815145121, 
    0.0448066281706536, 0.00263891698799167, 0.0329030526644576, 
    0.0175031548395292, 0.0257662707411015, -0.0321154304904144, 
    0.0187150890306518, -0.00463360681851051, -0.0194383676874365, 
    0.0489821021833648, 0.0990563680013752, 0.00137951557923642, 
    0.243570772269969, 0.255996312277805, 0.139666017973455, 
    0.0626085831895726, 0.120120301486325, 0.497178824966498, 
    -0.00166990380101709, 0.18219161266873, -0.417107123433129, 
    0.80362575627595, 0.3126463855506, 0.102668868994454, 
    -0.0945139585256387, 0.179714099840516, -0.119854198726627, 
    0.511979061645984, 1.06251273368631, 0.188820668508528, 
    -0.181177188124101, 0.128903668645634, 0.209101870080449, 
    -0.0814175365270873, -0.12892349924762, 0.0572076377435219, 
    0.0520338051196322, -0.0425650368901202, 0.0913157457960054, 
    -0.0349200282122054, -0.119915133940502, 0.0290265618214035, 
    -0.103392975951815, 0.0395212182927085, -0.11048175055817, 
    0.0491272369539194, -0.112429618124792, 0.0252992375170156, 
    -0.131757786619995, -0.0438464807654161, -0.00724643427670419, 
    0.0666936592486152, 0.00588404805673039, 0.0480944360059628, 
    0.00325756166923245, 0.0373040764572159, 0.0171866050512193, 
    0.0517282945643801, 0.0106427421606826, 0.0416851133089417, 
    0.0421302907236213, 0.0603621381910299, 0.0737043707490898, 
    0.0707459652771149, 0.0391614613141578, 0.0639480368928354, 
    0.0494157280727731, 0.0516868142616785, 0.0668602830816351, 
    0.0306904154971348, 0.0630635575145503, 0.0893940399482985, 
    0.144464798054419, 0.145028676437006, 0.0969034489707196, 
    0.103514939950902, 0.199272557001841, 0.161065186284764, 
    0.11273349676126, 0.0905592993500281, 0.0830870336317165, 
    -0.0728079296805768, 0.0546321864098859, -0.0541573606068341, 
    0.710100101067038, 0.443415962732384, 0.135572190267322, 
    1.10714680142184, 0.485084456161992, -0.0173725525412525, 
    -0.151323865353252, -0.0677160038148864, -0.107317852684526, 
    -0.0766287579193964, -0.070675494842344, -0.108289631485765, 
    -0.0503270491600355, -0.110165001228009, -0.0100677991086418, 
    -0.128664056797089, 0.0121313808222597, -0.0057965431170615, 
    -0.0114900885863976, 0.000627916811661008, 0.0498276241384264, 
    0.0318214188316961, 0.0810631081575039, 0.0799274269218044, 
    0.0535697303735175, -0.0570012899012072, 0.0387345747107399, 
    0.0926085375308903, 0.0963462708089829, 0.143928675315207, 
    0.184556002722239, 0.128223861062706, 0.074317316632931, 
    0.113150863932217, 0.178252943816046, 0.375865627039818, 
    0.225525374799447, -0.0898049869403379, -0.0782324627631198, 
    0.497700664524465, 0.370517004189957, 0.0901832329556137, 
    -0.214925293994625, -0.146464912939516, 0.420622736227859, 
    0.410640787218619, 0.106543315883279, -0.17582670955335, 
    -0.141700276150321, 0.417160880404584, 0.344852766491308, 
    0.104491886363213, 0.0584113525327283, -0.240166799289492, 
    0.490949786272942, 0.222982284736805, -0.119803383275582, 
    -0.0756852375163197, -0.148432110730814, 0.225216305482639, 
    0.0664839375388155, 0.0656565970372523, 0.162921530517613, 
    -0.0753159025853437, -0.0637244464478537, -0.111032430096799, 
    -0.284918041815566, -0.223534360864083, 0.0895526621799593, 
    -0.0931999003105398, 0.163716142999241, -0.0496907493099376, 
    0.154950981668917, -0.14975975492246, 0.107054880023389, 
    -0.213301358798198, 0.00320752455048259, 0.0688720743365176, 
    0.0649562447530995, 0.0874431921512515, 0.141951677416374, 
    0.109191547724994, 0.0738530635179549, 0.106380072114025, 
    0.0800589866817042, 0.0378278292511551, 0.132340315728619, 
    0.157642082207631, 0.125562741359132, 0.20934290876995, 
    0.266513763727987, 0.144447974576576, 0.12729863312807, 
    0.404857273059792, 0.21868478865846, -0.0994340604307145, 
    0.32873718409431, 0.444241271314489, 0.188217070813045, 
    0.133934175894822, -0.153761719305765, 0.435794164798693, 
    0.353246385065004, 0.129455614220744, 0.756890863641672, 
    0.543312263359687, 0.102750436938928, 0.0278208195881905, 
    -0.0169985983302217, -0.170900184762208, 0.118252406013697, 
    0.363215424640845, 0.136081177077602, 0.0620372662494079, 
    0.124139738780267, -0.166300430547749, -0.352014050474578, 
    0.00232618686715982, -0.253065782375647, -0.223732599472289, 
    0.226783402458747, -0.292311899940886, 0.0531247011320841, 
    -0.086902044872331, 0.0377127942836198, -0.26998953821374, 
    -0.00965845095138186, 0.112401677847622, 0.116270074847064, 
    0.159729025207143, 0.210350179463276, 0.165103693460894, 
    0.12183881967557, 0.161478124918927, 0.176817479629141, 
    0.147290507438444, 0.203521628752124, 0.186322682507142, 
    0.225134346069372, 0.380815629820663, 0.282605301290538, 
    0.0602846832185212, 0.179426565471971, 0.526407465125663, 
    0.326397507610163, 0.149763297953641,
  -0.0262496762553381, 0.417397070789579, 0.671233022739349, 
    0.17919027120702, -0.231976590020244, 0.105068366804754, 
    0.699390855924119, 0.0668086957364287, 0.167278325145675, 
    -0.261604889093158, -0.116062230513639, 0.417159997533036, 
    0.193256721032734, 0.0300778217939775, -0.0205645002377521, 
    0.0313457712168673, 0.000832496163716251, 0.104937331321782, 
    0.0772494543991638, -0.0156290575818063, -0.0466655986427334, 
    0.0415427170974423, -0.0749298789276618, 0.0081087790435735, 
    -0.123254909117536, -0.0673957990724186, 0.0245949971995277, 
    -0.0238702422979251, 0.129664008475501, -0.0521726989512118, 
    0.183574558937137, 0.0827207331135048, 0.0924728847942815, 
    0.44871043695136, 0.184643852579174, 0.0194987248908891, 
    0.0992901528325161, 0.373793372862576, 0.0886837839351888, 
    0.0695401498882485, 0.326790206165139, -0.0133031482106491, 
    0.241601135374078, 0.385188655304603, 0.27595138106851, 
    0.100640887626788, 1.17491268638512, 0.782410614862827, 
    -0.0293070900424307, -0.104312135826754, -0.16860185223757, 
    -0.185033500876981, 0.0927303242380152, -0.11165302733988, 
    0.119528737145796, -0.213828445568145, -0.00709473829949796, 
    -0.0394517867721847, 0.061712299895297, -0.208218685795407, 
    0.0105221413254697, 0.121767534836487, 0.123579521594845, 
    0.175767554179624, 0.282851965547578, 0.267218454005623, 
    0.200551392567025, 0.20118047006804, 0.257833934032825, 
    0.268687469719417, 0.260789746947654, 0.239323217947766, 
    0.20438617897176, 0.203699406711611, 0.287669567463274, 
    0.296223205766967, 0.172380138658153, 0.0531451055470571, 
    0.258476587116006, 0.412663461493168, 0.176807806480716, 
    -0.0426285487156107, -0.116387037011507, 0.275937077996116, 
    0.614837061553994, 0.332295401612891, -0.0712971928032803, 
    0.60670022665881, 0.251476978476471, -0.130571094700847, 
    0.228682508709425, 0.438454760373931, 0.249321830370199, 
    0.712611122924799, 0.185875852602644, -0.150248859490406, 
    -0.278707719506634, 0.165382553574756, 0.334126137635085, 
    -0.142327972857392, -0.11996200923209, -0.179681702199649, 
    0.0266656783579451, -0.198085874328247, 0.0266755017519907, 
    -0.170427342983607, 0.0200249440075386, -0.109219382990043, 
    0.0744354934379723, -0.186323994092649, 0.0391619542058741, 
    0.145435760422495, 0.151540543533621, 0.14933497406282, 
    0.204165979972035, 0.296503139828515, 0.347123275260341, 
    0.321817184846047, 0.255982710611945, 0.230217635208187, 
    0.33588012608502, 0.419707461726312, 0.371308386511995, 
    0.295699226611194, 0.330244825687549, 0.451900236688607, 
    0.427135912191337, 0.277573955330533, 0.209728142350795, 
    0.413026746799969, 0.468488715437784, 0.267094969171101, 
    0.142404127892572, 0.40019567150641, 0.437214217373577, 
    0.152815761607235, -0.0781810387180846, 0.238241798147512, 
    0.441851129125009, 0.277116918207712, 0.110208146428037, 
    0.00926404904513074, -0.321841776216542, 0.272662890870659, 
    0.482372700088298, 0.132355224225542, 0.102693555954325, 
    -0.090293769726449, 0.593003216405196, 0.00235676702841221, 
    -0.131528624452052, 0.0683038013149446, -0.00863678895017779, 
    0.148553027649667, 0.693842223981186, 0.112604721370876, 
    -0.027838238603015, 0.00359796830422714, 0.516492478264389, 
    -0.0589264838816579, -0.065860309780233, -0.1846842563899, 
    0.0957837667008355, -0.109815985269508, 0.0492157583366245, 
    -0.0783711446221359, 0.0924443204557696, -0.174298131691493, 
    0.0813074193416455, -0.257909240210149, -0.00787427960881481, 
    0.0307907849377726, 0.102267384440581, 0.207473062170547, 
    0.197751689277934, 0.141558859887409, 0.117539144598397, 
    0.136679464630075, 0.164863046921481, 0.252202519143996, 
    0.27205985169217, 0.0556502648964278, 0.119089884588892, 
    0.621955047407453, 0.265088754834666, -0.0873249426815097, 
    0.297129205230276, 0.50969420810923, 0.139436705834844, 
    0.115389605757533, 0.0947098945231119, -0.0244957452409837, 
    -0.344532379211509, 0.847768397379556, 0.212143949257379, 
    0.0775863620713117, 0.0387184161359993, 0.0737015683689416, 
    0.141857194944406, 0.0300367801744896, 0.0149904031494484, 
    0.530552393383438, 0.447592402818638, 0.257214397371648, 
    0.311575112636472, 0.328680826436395, 0.155226914218259, 
    0.0416614805770983, 0.065389847350939, 0.225676007649987, 
    0.216351704747199, 0.12292711474842, 0.117726675637475, 
    0.239928032187486, 0.220539828485248, 0.109402773951818, 
    0.0877072271439728, 0.186551366312733, 0.0802303209575028, 
    -0.00521954719124253, 0.594500069427401, 0.158041549630325, 
    0.00699573068700871, -0.134643628262538, 0.453963756754436, 
    0.414864955770782, 0.195725831276716, -0.131336998605327, 
    -0.0274127247505522, 0.401505436131927, 0.479022178720713, 
    0.173819367618333, -0.225692700190332, 0.13663959133452, 
    0.438453414943884, 0.366133180181872, 0.248320149861229, 
    0.00652004167178055, 0.697278953900745, 0.210813455023048, 
    -0.0340904045827531, 0.0944749731517742, 0.271018242122199, 
    0.0346193737950327, 0.158243742310564, 0.430109474366425, 
    0.308949347611404, 0.15603060518394, 0.325229360128473, 
    0.385178204251878, -0.0220001550900735, -0.0537595848469523, 
    0.0510420621096013, 0.068199401298491, 0.0298272091426658, 
    -0.0117701630953954, -0.0798063274334518, -0.00152893956547555, 
    0.0351766175545482, -0.0462642391087817, 0.0191466623179615, 
    -0.0436842700205874, 0.0444743782580041, -0.018418182691278, 
    0.0407038770835349, -0.034956781944668, 0.0391403539333152, 
    0.000153426777126875, 0.0750650152576195, -0.0393061899863212, 
    0.0953575964450968, 0.0211640486642964, 0.36451495928169, 
    0.228571831876233, 0.064548048944675, 0.162628742447633, 
    0.262572374802424, -0.0471672774580896, 0.335794420124478, 
    0.512972680692824, 0.0736059650845542, -0.0823109519311501, 
    -0.365728547308266, 0.451889607448383, 0.5031186585403, 
    0.701301445632767, 0.462022449486252, -0.383905879315837, 
    0.437135137413368, 0.6520784944819, -0.142512776206438, 
    -0.132946949071591, -0.209434397135968, -0.217797116606554, 
    -0.0849836515441776, -0.105058072307754, -0.117220652092537, 
    -0.272107921940826, -0.233543121446593, -0.0303384465032801, 
    -0.0801659950430095, -0.032265004723313, -0.252960507266696, 
    -0.0550887196194755, -0.0363441481114338, -0.263400401126252, 
    0.0254649987304096, 0.0266999650024918, 0.0340418278262585, 
    -0.207913130400661, -0.00850377387085317, 0.013589345253506, 
    0.000617903041592885, 0.0643459113776351, 0.0275630904989823, 
    -0.0215312711941956, 0.152229278187936, 0.0501783637364015, 
    -0.0455286183606223, -0.224725301577531, 0.220706810838888, 
    0.123038351938415, -0.320762601569604, 0.667262342363811, 
    0.42063736825252, 0.108296214921735, 0.0798142806655099, 
    0.308071402494787, -0.231037100386536, 0.588966893529178, 
    0.391529050099499, -0.0170727253884239, -0.0542702492365419, 
    -0.0391291902121421, -0.025568532282232, 0.00644167506521533, 
    0.0323164419880655, 0.119492261778625, 0.0133510365018551, 
    -0.0188645885656845, 0.00132912319534621, -0.099216692308839, 
    0.0832043788968457, -0.0863314125250336, 0.0579773601590685, 
    -0.0966559564796684, 0.0576895515572719, -0.126953166024871, 
    0.0279368539540238, -0.182160238985599, -0.0475463487066822, 
    0.0368703989970364, 0.00331516945803849, 0.109391797579243, 
    0.0825200295059944, 0.0150966385196342, 0.156904727908673, 
    0.115147271175544, 0.103958860597081, -0.358680985381622,
  -0.284434250099961, -0.0936070916279582, -0.298496384512662, 
    -0.219828950570702, 0.193138123252716, -0.400494500289413, 
    -0.0140354239057261, -0.112318503447777, -0.0396860051396868, 
    -0.262946108028835, -0.0479371342300679, 0.0284555318228161, 
    0.110140432177662, 0.130125644209409, 0.0995933438217606, 
    0.0696893126367953, 0.0972836132257375, 0.160187088282301, 
    0.12443683638845, 0.0628785601054223, 0.135381059980175, 
    0.20866692072961, 0.202631797428313, 0.143648907510414, 
    0.196551390909512, 0.311463922030956, 0.198106634146654, 
    0.0249760371171127, 0.174329108713324, 0.446916049382991, 
    0.109020957552951, 0.00901282225704485, -0.312392091778952, 
    0.260021151230664, 0.380702298582759, 0.719158290941472, 
    0.373270225928347, -0.1408765200423, 0.0701761491939721, 
    0.630216667519558, 0.242615288645832, -0.0494986897785842, 
    0.695527777811811, 0.363099835475499, -0.105910290897671, 
    0.888768322640171, 0.44418743668098, 0.00256204098173604, 
    1.00418998252247, 0.483623797147053, 0.00938354638300027, 
    0.00716377874594157, 0.00344750775080099, 0.00439265910193225, 
    0.00863807821139677, 0.0222647868361957, -0.00626918510696499, 
    0.0532362942572777, -0.010375709062266, 0.0644816054579229, 
    0.241113097766525, -0.0686143462131097, -0.147754601562347, 
    0.319680521947972, 0.434913094554406, 0.22151886831865, 
    0.195294385533982, 0.611251963788856, 0.140786551391179, 
    0.238004215146606, -0.57497352453388, 0.331953299480156, 
    0.557719565848292, 0.207118638104547, 0.123510153380578, 
    0.134243939416596, -0.371658449485004, 0.43776038435138, 
    0.670505212631065, -0.43227220238534, -0.195991217611255, 
    -0.246466023626999, 0.03526945815184, -0.167277027010694, 
    0.0637465420562146, -0.208954765288956, 0.0492979994560084, 
    -0.258705355947943, -0.0073761159567723, -0.165442003797739, 
    0.0578354528821113, 0.0449649362005932, 0.152790074977248, 
    0.215426401208115, 0.225147051636116, 0.28355505646214, 
    0.249498541153661, 0.136734147199188, 0.148942569576439, 
    0.28194492696362, 0.201902887122708, 0.142297182891893, 
    0.129371885051344, 0.125572129213088, 0.116416527954447, 
    0.134417928020096, 0.141176304817173, 0.126385411839221, 
    0.126251124557378, 0.13704740344538, 0.113259587569602, 
    0.0950621964445389, 0.100062458746555, 0.102180279390389, 
    0.118543740020413, 0.0934842415899572, 0.0564500951528269, 
    0.130829427623362, 0.123770766860595, 0.0445276786687217, 
    0.0567018227278222, 0.0336660091584159, 0.546667299368134, 
    0.299091152055746, -0.0704598783542421, 0.276357328298861, 
    0.536444296811812, 0.227699703730424, -0.101886386942096, 
    0.244089225072574, 0.611742906363158, 0.612121662485134, 
    0.486070372081104, -0.46377688365314, 0.239091779683173, 
    0.570437694807228, 0.329530182731075, 0.225435548885968, 
    0.0548799411346205, 0.539933030308752, 0.574426167995069, 
    -0.0216186268045406, -0.0969666269531877, -0.162124217996426, 
    0.117696046111371, -0.121553192032732, -0.0749933764409079, 
    -0.0912796974982761, 0.0632879279782924, -0.0333398876598586, 
    0.0520523526525207, 0.0360850386069743, 0.0911615001266825, 
    0.0788531259037387, 0.0674094153499974, 0.00180710649339057, 
    0.0924268312305343, 0.0936980283692278, 0.0511236527795552, 
    0.0084060536309622, 0.0673317575107513, 0.134370279853329, 
    0.124476659809869, 0.0885422299760857, 0.0804030434117172, 
    0.114028022827211, 0.107390964658485, 0.106227788686254, 
    0.129656063469979, 0.113783980806587, 0.0631443225450219, 
    0.0457914421352773, 0.0662272935442807, 0.0682864257612967, 
    0.0748557557060956, 0.047183519242075, 0.0611883963131875, 
    0.0878025390887319, 0.085661136472054, 0.000690774921928941, 
    0.0671821615206616, 0.214779638524945, 0.153303038442533, 
    0.0450919475231914, 0.194705971249997, 0.241513725490358, 
    0.165022161895359, 0.359145451060145, 0.297181294156738, 
    -0.0202015038622162, 0.640875466007618, 0.331773212077604, 
    0.0331765711847964, -0.0914259040904143, 0.403884639287944, 
    0.575928430159019, 0.355418873584338, -0.00086065277524186, 
    0.541028046050414, 0.245804355331442, -0.0660553212454623, 
    -0.038514499598907, -0.0409057097777658, 0.122521471765348, 
    -0.0464295442455497, 0.172731942418561, 0.283370034927014, 
    0.0686740561133892, 0.131681363810907, 0.186462411650104, 
    -0.0791599727532612, 0.13194600133085, -0.121913650084824, 
    0.0845240779021193, -0.160216661866026, -0.00704727317350212, 
    -0.343103752600303, -0.148397574989773, 0.00536102260964738, 
    -0.273797450791946, -0.00116741513812961, 0.066277556121873, 
    0.0761844898038974, 0.0916186564516863, 0.111489773271597, 
    0.0958164489343732, 0.102132481189854, 0.150919095637771, 
    0.106608648235776, -0.0185743396387343, 0.224793243629928, 
    0.256627709731597, 0.0609512234397519, 0.0891450174516453, 
    0.440723262900608, 0.274512432411033, 0.0834418456818993, 
    -0.0719617498344899, 0.1492362675695, 0.577500897307622, 
    0.170819276031155, -0.0311368781834788, -0.0815012881808906, 
    0.232617351100936, 0.169844165133254, 0.534429433812125, 
    0.516732857037256, 0.0475054119646731, 0.486697342729812, 
    0.6980475229277, -0.158685298975507, -0.098878304331541, 
    -0.0799645570873302, -0.103486791967301, -0.0366438126338108, 
    -0.105823561267892, -0.0505614324779967, -0.118810556565765, 
    -0.171840559794224, -0.0516801960799412, -0.209863034880372, 
    -0.0533546095546077, -0.0345709421251012, -0.146078828763868, 
    -0.0574042190011891, 0.0278488543526953, 0.0302674309623626, 
    -0.0106947864864972, 0.0963902869609276, -0.153211058764114, 
    0.0176720654156252, 0.0387443039991137, 0.0625718157798398, 
    0.0942083515560147, 0.0995146683587659, 0.0836713182373221, 
    0.0916898006156196, 0.150420872698454, 0.106201677014152, 
    -0.118628942216577, 0.227075924944863, 0.382182451894064, 
    0.126530466359111, -0.158577454017667, 0.105742087496728, 
    0.450483906561284, 0.396896589973291, 0.186419368184951, 
    -0.262774036790849, 0.219975004838091, 0.440877035482919, 
    0.12054635049875, 0.242170626889338, 0.570142649583249, 
    0.387288772890723, 0.104818242126774, -0.316770873861635, 
    -0.223432229915599, 0.535624948354501, 0.220257656034941, 
    -0.043668995839434, -0.012696445422734, -0.12362678443903, 
    -0.0917012031770649, -0.118445721999005, -0.0733688415824504, 
    -0.0973648749467602, -0.208276940977121, -0.0430390105248387, 
    -0.138418228116886, 0.0414358797570746, -0.126792793775568, 
    0.0218487126420077, -0.061655752223027, 0.034003786972345, 
    -0.0842246987703938, 0.0324698585664333, -0.0264117721784558, 
    0.0728372902089831, -0.107779703672722, 0.0577383354350592, 
    0.0553890513029448, 0.0554657209743002, 0.0536981254390094, 
    0.0581085711502241, 0.0599874588784563, 0.0683162373526402, 
    0.0756679058775283, 0.0647191811058324, -0.000304867173867795, 
    0.115117390539824, 0.172992606797328, 0.103569481991361, 
    0.115910529993851, 0.280327907963744, 0.172971885060336, 
    0.193760313732854, 0.38732548638892, 0.113631992445088, 
    0.0564979128810383, 0.250584607780877, -0.294574017800589, 
    0.420426963848835, 0.409921301763104, 0.170151402233735, 
    0.379192107318643, 0.429020451243007, -0.247676235333408, 
    0.504158336415857, 0.464555925828454, -0.220624042831433, 
    -0.14392840357809, 0.0438652873389535, -0.179553833857787, 
    0.0390087915986688, -0.0897541281376082, -0.131699929990054, 
    0.0506935478143664, -0.140459873615226, -0.0823835615845037,
  0.341700677875003, -0.000826372939201542, -0.065101077606427, 
    -0.0652079326147593, -0.0603157526352467, -0.0612153434295116, 
    -0.13815763508027, 0.0900392146322936, -0.101858539750541, 
    -0.215406248586891, -0.0979249898884571, -0.128480054590231, 
    0.00059895363219109, -0.144921021605153, 0.0479956696596415, 
    -0.139002734705623, 0.0563768370365757, -0.0658659556842459, 
    0.107375301511744, -0.118140346554781, 0.0670081252459312, 
    0.0232382930639943, 0.0525624464219338, 0.0321733025401279, 
    0.0515232833943962, 0.0135665440577064, 0.0360274824492724, 
    0.031660385141357, 0.0443452579592403, -0.0129879249920044, 
    0.0419753815865733, 0.0738613134305998, 0.0802260321942966, 
    0.0733073815127552, 0.0792304295418508, 0.0661932919746977, 
    0.0715759596160608, 0.0739852295933882, 0.0723679259077392, 
    0.0235030633999812, 0.114965121445379, 0.14867680012685, 
    0.0959775768664889, 0.122096851598523, 0.277298065749817, 
    0.214838872500453, 0.0829469019408086, 0.0314281342476732, 
    0.224537062447385, 0.301050891358403, 0.270065323699106, 
    0.100568427281773, -0.0116413947870751, -0.200324014428222, 
    0.543072421274556, 0.359059805123946, 0.0638871821364334, 
    -0.0152727767897046, -0.0157945358072442, 0.562537963336002, 
    -0.0437674745269359, -0.0584552324860628, 0.0173936391820383, 
    0.0714960013330626, 0.0421546565740623, 0.309830634188535, 
    0.0977935871579381, -0.136351315704308, -0.1894790860981, 
    -0.0827058832774673, -0.246799939516197, -0.421588555762842, 
    0.347295311732207, -0.149633662651309, 0.160086120340711, 
    -0.374624424910265, -0.0729430297411315, -0.144078973373663, 
    0.00703669963462354, -0.36015583299644, -0.0430046391956913, 
    0.149762473474414, 0.0612320004057979, 0.153119572546044, 
    0.386760040983146, 0.256624002944062, 0.0850181030351302, 
    0.1388277803705, 0.399911797196739, 0.257944124764061, 
    0.0781348640753311, 0.0283458337043845, 0.117046132666499, 
    0.0665946407454633, 0.0891214557229866, 0.0661353251125249, 
    0.0662237601677291, 0.144251660306405, 0.133596458979919, 
    0.0251992084581091, 0.116513555222529, 0.213826190213754, 
    0.0466943197684596, 0.1118838316245, 0.264553043542834, 0.41850239505223, 
    0.256473976925679, 0.0240154459545443, 0.338699650994773, 
    0.260731546900167, 0.13726488668416, -0.135886076861799, 
    0.756675874930056, 0.490830470960573, -0.248576832712682, 
    -0.0443349930520661, -0.63967064999215, 1.16635625451723, 
    0.0579188688011308, 0.0284593198377636, -0.233570371464216, 
    -0.0864019023660239, -0.0246096261868551, 0.064760553288673, 
    -0.0993109532655268, 0.044854162929615, 0.134561049141215, 
    0.0175265750659701, -0.0191941438864842, -0.0267153593151861, 
    0.0383550030969886, 0.106709137265759, 0.0155539684778773, 
    -0.0151011359256896, 0.0339584622134042, 0.0132365092737282, 
    -0.0256381823773691, -0.00469961544965307, 0.0113093224575721, 
    -0.0790442886275468, -0.0333797992332891, 0.00182051198051263, 
    0.138451765627812, 0.282456436781081, 0.304016480593698, 
    0.20644547574948, 0.0931067466816815, 0.0103703939050601, 
    -0.0706285933143494, 0.265753015855039, 0.4320239148342, 
    0.205230247832703, 0.113590681933205, 0.502479549751511, 
    0.30979772013955, 0.0328895138297877, -0.0916874835531415, 
    0.517786438487552, 0.426925219603545, 0.182279826299574, 
    -0.142270710036679, 0.351213744452185, 0.399358763993517, 
    0.152475428631115, -0.0951361816840466, 0.273846758446103, 
    0.256538717090515, 0.121148412734367, 0.599368491982133, 
    0.356947327311853, 0.0355695234939839, -0.0596121333440557, 
    0.424263086472365, 0.141103407003642, -0.0208703170032976, 
    0.0371440201754562, 0.332389633043395, 0.168541369802171, 
    0.0457727011116465, 0.0465088566219295, 0.179213744947722, 
    0.205229361205032, 0.170426578883782, 0.196234300453177, 
    0.196096592094696, 0.111889120509532, 0.0565518691897964, 
    0.188235091171968, 0.270885834905661, 0.136606129714834, 
    -0.110279694168914, 0.157855583878814, 0.404309866056682, 
    0.156270097268987, -0.0464744089818119, 0.155844331018222, 
    0.486257994429471, 0.383120076909022, 0.116285272505244, 
    -0.401650228324062, 0.130569302204091, 0.488622498265884, 
    -0.0789389259668015, -0.159347489274107, 0.15366729251125, 
    -0.023448346858213, -0.0143986407826958, 0.705841957482875, 
    0.216652531876715, 0.0091560339577799, -0.195691443311636, 
    0.0773972142974443, -0.16248893429791, 0.0041379611111993, 
    -0.26792237398597, -0.0953905611860044, -0.00337152363857035, 
    -0.0861421596758746, 0.195671232417803, -0.204831940665473, 
    0.00981001233166972, 0.165178817189325, 0.135565161463386, 
    0.0584901685979468, 0.117819514945481, 0.294680489583803, 
    0.338803085519404, 0.266779497467778, 0.163307407695942, 
    0.121393219986933, 0.345531934268399, 0.312582845722144, 
    0.193278948529983, 0.529296481440186, 0.559908502760555, 
    0.193012732409784, 0.0301384743197862, 0.731054776588254, 
    0.383749191498598, 0.0322868459595187, 0.039751034081635, 
    0.736562110533617, 0.111611328440558, -0.225898134410721, 
    0.182023630142771, 0.528133196945581, 0.153083021309283, 
    0.153392399404357, -0.254929884621028, 0.309897812053372, 
    0.331061980572489, 0.0523776159412504, -0.0224823981470769, 
    -0.0766241790312217, -0.0160279174058723, 0.0484410086836748, 
    0.756735365748918, 0.269180855803961, 0.0716954361672356, 
    -0.0017891199664161, -0.381780148825846, -0.158293599242099, 
    -0.102318718691444, -0.272314071429936, -0.0477772478041596, 
    -0.278626302508877, -0.178221872434005, -0.0412117299229688, 
    -0.240179032487905, -0.0375212024548949, -0.0778365978937476, 
    -0.0195753350177872, 0.0301599974287562, 0.0232615146734941, 
    0.0990793600477769, 0.0522273302904724, 0.0772018150979798, 
    -0.00915009339892992, 0.0567994673777977, 0.0236612510631997, 
    0.0736310199945949, 0.00856336611586434, -0.0284447912273292, 
    0.0486142720172014, 0.0889640563001323, 0.0907343252824149, 
    -0.168304056546032, 0.219226804063699, 0.204108175336831, 
    -0.195063662391874, 0.222778451764738, 0.114277870496192, 
    -0.390423790418061, 1.07703147265905, 0.63605579753733, 
    0.0530077429795546, -0.488021641322323, -0.0654583879656095, 
    0.743033762319542, 0.428109884931176, 0.166645226012989, 
    0.286276232890763, 0.203601753297587, 0.112221147512089, 
    0.113011980261732, 0.129431603688978, 0.0663748203104262, 
    -0.02897690381778, 0.131146630606094, 0.110310104975091, 
    -0.0440060043163114, -0.0413510837720607, -0.0589549155163819, 
    -0.0572879903561637, -0.0292347146101325, -0.0668625602595219, 
    -0.0315247190349352, -0.0379354448280084, 0.0168007283781358, 
    -0.106260999936718, 0.0634664767291265, 0.171208346310844, 
    0.116707397372646, 0.0232518802073849, 0.119331677238669, 
    0.29717329009766, 0.205894814852351, 0.0906996493590381, 
    0.0645121633174223, 0.200358218795047, 0.277286398451061, 
    0.213212442759534, 0.15899445171741, 0.194773410448389, 
    0.251776987323001, 0.188771961500977, 0.0984787971063749, 
    0.17797280657287, 0.339235378506385, 0.174892182570812, 
    -0.0490115081518138, 0.24436089729416, 0.420590567877228, 
    0.133638248026912, -0.146566156794309, 0.415387600664108, 
    0.470184957722251, 0.021853953003088, -0.0450730117765474, 
    -0.274142655539512, 0.471570154769864, 0.366585085594348, 
    0.126205944782678, -0.0288282301342357, 0.0709148544265676, 
    -0.23180908752076, 0.52081406833946, 0.518211516364737, 
    0.183423260508335, 0.215082936099203,
  0.47740194153648, 0.00822538967437938, 0.0968090422438452, 
    -0.337223278521818, 0.22046253657245, 0.43361779970475, 
    0.269221284190155, 0.177196723000503, 0.13693544889877, 
    -0.157413831809674, 0.197325803013154, 0.438487270346544, 
    0.142699956985153, 0.0310857545835224, 0.25263040150919, 
    0.129987851715102, 0.145036270364146, 0.506974427046436, 
    0.195988328700151, -0.0132607573249562, -0.0633645672607156, 
    -0.235557157855917, 0.0951227365239142, -0.121794544063349, 
    0.0771639221820216, -0.220413701042972, 0.0607733307891891, 
    -0.368411068945151, -0.089245682591654, -0.150201659590411, 
    -0.105456787773071, -0.0190276029205366, 0.131098976380292, 
    -0.0137711842207375, 0.121657178551298, 0.163490042322313, 
    0.071245249224919, -0.226068417420587, 0.116493016700441, 
    0.271098523327961, 0.149208842782282, -0.156750016285965, 
    -0.193706918766935, 0.687412639092238, 0.471673386567244, 
    0.349474179224705, -0.452330812683919, 0.749963936947093, 
    0.600663699824948, 0.186050249930523, -0.0965877867643334, 
    0.143761252188562, -0.128202495368307, 0.010072705220108, 
    -0.0525491058671186, -0.0548537428330524, 0.00846386011901299, 
    -0.149411864070569, 0.063636045904803, -0.048986102196278, 
    0.137149452640689, -0.117193759541337, 0.0494939244103915, 
    -0.144952645587989, -0.0891686949382337, 0.0213267843784588, 
    0.0702714313042617, 0.0214890846525376, 0.115227370468464, 
    -0.229080636296515, 0.0345657004802498, -0.049512587834712, 
    -0.0429809187414151, -0.0150228055982669, 0.0276339371600552, 
    -0.0278221360871677, 0.0208215180209948, -0.0111539117796821, 
    0.0208166694774258, -0.0803357490100042, 0.0218073156606213, 
    0.0756376539476654, 0.0765987697417647, 0.109759096891128, 
    0.1576447969407, 0.0920976147678992, 0.0220870275512754, 
    0.395401018433212, 0.0781279589474226, -0.290158766089625, 
    0.0784340194976466, 0.470613762555575, 0.0405102289782464, 
    0.468020081637033, 0.566260456365072, 0.281038832845066, 
    0.297540412351835, -0.312876431759099, 0.379362413227263, 
    0.454834187036454, 0.0524346717790137, -0.0386254098005047, 
    -0.251739616871219, 0.601498074253356, 0.220816775382649, 
    -0.0365506553692249, 0.0277375719001012, 0.250535671792603, 
    0.395787929802284, 0.507181064719455, 0.232496166509879, 
    0.0229159911424952, -0.0356831841660474, -0.0620843353704272, 
    -0.0725008495054654, -0.0937817981395247, -0.109999339364026, 
    0.0670830445824348, 0.0697732078792735, -0.162935154430034, 
    -0.169277025177211, -0.0627920558170077, -0.122899042563296, 
    -0.0339257094533362, -0.126296495122511, -0.0524340596949778, 
    -0.0959252329358218, -0.0719299126464461, -0.0815377376415687, 
    -0.0392540055118542, -0.07459365373931, 0.0254776313316926, 
    -0.0933558123496165, -0.00830736736697604, -0.0174185262575817, 
    0.0485145069903807, -0.0889033875272057, 0.0113530904222591, 
    -0.159016749807062, -0.107306659873565, 0.0310780885103647, 
    0.0415447511328146, 0.0635535145092243, 0.112361518613039, 
    0.125645761482431, 0.107466405908255, 0.0994760079307251, 
    0.109253543365506, 0.0851842387170627, 0.116869529731888, 
    0.255563765944792, 0.114841421435262, -0.0356996584214136, 
    0.0322043482206105, 0.555186328485092, 0.382558097488551, 
    0.0805598996225953, -0.153433068238205, 0.11987129268277, 
    0.365844817421865, 0.0434707769513598, 0.992282979703839, 
    0.443805692268999, -0.190458605641257, -0.067041851265285, 
    -0.0486003455014468, 0.671588308660437, 0.0149535086530591, 
    0.899210150556531, 0.77576885438026, 0.00878094559479332, 
    -0.00435414766081636, 0.00953404427885814, -0.00903471094641863, 
    -0.00121101303367353, -0.00197126449000139, -0.00039435273830743, 
    0.0101662995749425, 0.0164818287459172, -0.0365200996058266, 
    0.0284446855390568, 0.11913410927894, 0.16428814239347, 
    0.130166884460723, 0.138110733674731, 0.217905741054313, 
    0.225666560600777, 0.161830533746174, 0.101846052784698, 
    0.0904375763587199, 0.226185343302788, 0.267812251427116, 
    0.209241011908816, 0.196962746553586, 0.258176151662364, 
    0.300353741518636, 0.302037890100893, 0.183039445940142, 
    -0.0296459922484816, 0.15361167602395, 0.53789259436432, 
    0.199183351935357, 0.0386637591991854, 0.000675362478436539, 
    -0.137428568533872, 0.664344168833194, 0.275168106121462, 
    -0.0505374861763694, 0.321341891737555, 0.407272661492843, 
    0.0648556576165003, 0.532625306604992, 0.302051963103805, 
    -0.223340584699986, -0.0686977647988068, -0.113368479539608, 
    0.510727948470091, 0.142041324108434, -0.172255522417686, 
    0.516153426663343, 0.266914474758208, 0.0799501907986751, 
    0.0422554916738013, 0.044034477856961, 0.0604400283329372, 
    0.0449179113072079, -0.0145427737345222, 0.133897097824582, 
    0.113220865470033, -0.0539481215720246, 0.118184816480081, 
    -0.00623036478872631, 0.230842205326361, 0.50595009035071, 
    0.22546478355053, 0.0912228017411698, 0.0759095229530934, 
    0.120882080238571, -0.206097241819594, 0.189493301583351, 
    0.646431267832733, -0.0422655738866426, 0.0217569028109417, 
    -0.340989007946609, 0.295666519106237, 0.534527946872962, 
    0.369722351969279, 0.139513304703098, -0.175564352117282, 
    -0.0513685950608497, 0.462306418753145, 0.268369055619276, 
    0.0847857296295166, 0.0429833565291891, -0.0732560002716487, 
    0.0847362758319257, 0.0815529556304914, -0.000231699990481865, 
    -0.0153770788698393, -0.109070697871471, 0.159179681962302, 
    0.192093627651012, 0.0904317599808358, -0.00245456441947725, 
    0.0836330466886893, 0.223876264227874, 0.213997166622341, 
    0.126743565632464, 0.0397740165011175, -0.21118771676918, 
    -0.00381716835318148, 0.541596305775912, 0.151862330531605, 
    -0.00127657244241641, -0.11161853183816, 0.535501643244006, 
    0.200623299096683, 0.0286896604498214, -0.0724100438565019, 
    0.439937740692913, 0.270413241406372, 0.0898902503770352, 
    0.0190848959909034, -0.0469671348430426, -0.00325515108312917, 
    0.124544956015656, 0.392093235090738, 0.0782311165896915, 
    -0.0735198673860665, -0.00813724246116317, -0.179716173349489, 
    -0.121997051671108, -0.0728617617512397, -0.153620597668839, 
    0.0193718199662846, -0.146844090029262, 0.0274652450720854, 
    -0.0637056885063814, 0.0745519324003223, -0.15716765940894, 
    0.0142946171531497, 0.104279678532786, 0.136270143076682, 
    0.141090575083865, 0.149650421616166, 0.166166266423975, 
    0.15708903490394, 0.143013962380327, 0.179509587740556, 
    0.186755769238619, 0.159230037442735, 0.165230394225987, 
    0.158382941779425, 0.118089484895642, 0.134319977127276, 
    0.124783807987023, 0.0955996727824914, 0.0667414091026098, 
    0.00289139169852295, 0.132857698793993, 0.266563229989323, 
    0.177640459907699, 0.736199510077472, 0.300111499711935, 
    -0.301043757815052, 0.417980865111234, 0.444160384257445, 
    -0.22469068657534, -0.126874344057125, -0.0135894232902107, 
    0.264668492682848, 0.0763418125257125, 0.00970511580614369, 
    0.0121903659977246, 0.123557818106517, 0.0555226150800531, 
    0.0915965993194105, 0.190983138782116, -0.00657624982745234, 
    -0.0582539576548798, -0.0403744004562375, -0.151090625918224, 
    0.0652734663941223, -0.133463346529635, 0.0371403190295868, 
    -0.138149243005112, 0.0233639863674545, -0.273892129662633, 
    -0.0695140139473755, -0.0945556624129275, -0.179247636045195, 
    0.0205975103212574, -0.144173827384802, 0.00350888221903124, 
    -0.196969473199254, -0.00815532221835376, -0.192972906244475, 
    -0.0992239426056792, 0.108688821199512, -0.102571835332653,
  0.208315229696631, 0.10999666895016, 0.152458320848993, 0.568559828585137, 
    0.0548300386647356, 0.00676459590858396, 0.0376666335889894, 
    0.415553703614901, 0.0514680285062942, 0.00708875265744136, 
    -0.138096725118697, 0.284218282511783, 0.275483881171992, 
    0.114113155851401, 0.0506552507294789, 0.284925677059656, 
    0.214432953255007, 0.023052900320321, 0.0520450036855483, 
    0.405297103392474, 0.253557604606823, 0.0887309161684408, 
    0.0766155823712552, 0.271620724751082, 0.237122261764424, 
    0.140852400428435, 0.132159360619479, 0.210372252838314, 
    0.437146649709014, 0.24501216212546, -0.0670269247951995, 
    0.248842902592602, 0.396293030231861, 0.240422895412576, 
    0.399275877427823, 0.350841987320223, -0.232380245500071, 
    0.452680924232502, 0.56860606134035, -0.135440752051998, 
    -0.292145796708131, -0.0677126290058185, 0.400699339832007, 
    0.144924564971028, 0.272826325048545, 0.548866748679664, 
    0.140727986647767, 0.123154289167258, 0.774554654189975, 
    0.17065309523461, -0.0363517631802683, -0.00569385293282156, 
    -0.0355864862451498, -0.0111396239014055, -0.0348822137255064, 
    -0.0156352566550422, -0.0294053163336121, 0.0333070455854318, 
    0.097327083103621, -0.126390627222617, 0.117075758841795, 
    0.226609307064303, 0.00618408085677663, 0.400428647915311, 
    0.315938007433483, 0.133888830294693, 0.503886819273977, 
    0.274734200130661, -0.0634749789093361, 0.037154238612403, 
    0.682461167282957, -0.139503767459024, -0.401880062136752, 
    -0.175732173922203, 0.983878040799383, 0.170182296908171, 
    0.0323133020996395, 0.443172580160024, -0.242250982432021, 
    -0.30287197465802, -0.115786162539415, -0.289761611538571, 
    0.0042753505558579, -0.300546084392389, 0.0966369021396366, 
    -0.394275830869269, 0.0249027038710988, -0.375659138587065, 
    -0.125505909124921, -0.21619918248279, -0.083371630945322, 
    -0.0161160356002573, 0.0411269156244068, -0.129330158118906, 
    0.152680031888251, 0.0692099636811319, 0.117726271548488, 
    -0.00688683712401253, 0.0384510001296968, -0.163889620568749, 
    -0.038466752295066, 0.00944599360425224, 0.0118443979089073, 
    -0.0344938077946419, 0.0772074024149769, 0.0765346083100651, 
    0.0549337469857545, 0.135858224994369, -0.0826502289173995, 
    -0.0754222947211354, 0.391310872491043, -0.163598375820301, 
    0.341662516068983, 0.472430197524283, 0.41805830949525, 
    0.250941868309101, -0.0361897037779848, -0.0247307605318278, 
    0.633874828157178, 0.219933745192659, -0.080289905915001, 
    0.724720707292918, 0.442043602970961, 0.134648927495336, 
    0.179000196850271, 0.430685989054806, 0.241747755518571, 
    -0.121840523660574, -0.351054982480293, -0.146924010645035, 
    -0.252623023693641, -0.224576423657873, -0.284606692400058, 
    -0.0811047484719443, -0.268918087194003, 0.0403130869241079, 
    -0.203779803285515, 0.0422123830127378, -0.339625906420613, 
    -0.153187986272647, 0.0288517229593445, 0.0885588270200067, 
    -0.0330515829446681, 0.0120730310836204, 0.0854110190053763, 
    0.0208948834560147, 0.0888473972709167, 0.0876569984840268, 
    0.0992939431095057, 0.0341683061631842, 0.0424477931283711, 
    -0.0138900438017932, 0.0099891887570438, 0.0128500031320668, 
    0.0223622821755209, 0.0135886237612211, 0.0303112155351323, 
    0.00718844227175679, 0.0459544743625662, -0.0230756486068865, 
    0.0469848540037888, 0.0822027406852394, 0.090331610820913, 
    0.127560731063077, 0.135969408316415, 0.067281323840661, 
    0.139364316927212, 0.279983849193181, 0.0104476254976122, 
    -0.00808339609087772, -0.294183696221741, 0.251376275170237, 
    0.452077243944192, 0.161998950850985, 0.0256452689059986, 
    0.00537792103883612, 0.0676402374728524, -0.00441812865251603, 
    0.649850141893526, 0.507956975818573, 0.0995809596176539, 
    0.0551355572064923, -0.0929317958523702, 0.36988253114812, 
    0.273903247975759, -0.0221857102811077, -0.0950680710381678, 
    0.565855270557338, 0.296167983888966, 0.0317924684707089, 
    -0.167214284814769, 0.107976718393288, -0.118386296438135, 
    0.0744087796017353, -0.12658311887391, 0.0517071783249611, 
    -0.273236463467425, -0.0564061564169738, -0.30721863984792, 
    -0.239625941413131, 0.0318730081506923, 0.0243388393997564, 
    0.0646693600928866, 0.0338694403428444, 0.0416938462852142, 
    0.0614945452849063, 0.0827101172606128, 0.0751030422206448, 
    0.0854314552302865, -0.00850394861275432, 0.153132683271713, 
    0.184183716441181, 0.196982268615382, 0.252786849528933, 
    0.135219600869315, 0.135841991565138, 0.456550317130464, 
    0.18259039285728, 0.0690873457150238, -0.189748727437691, 
    0.483956753987779, 0.460713180205649, 0.31970030462391, 
    -0.183840035859963, 1.02276178491695, 0.692318430272592, 
    0.415805647657998, 0.882900728441239, 0.11715862584923, 
    -0.221409660278477, -0.135793866759411, -0.191448731156737, 
    -0.199490973611891, 0.0559873140039156, -0.119600474209245, 
    -0.0241864012960179, -0.0731014612135265, -0.157062902007335, 
    -0.044695522634242, -0.0706848664668093, -0.260198108617574, 
    -0.00630465815231837, -0.027275111692778, 0.00392369246851806, 
    -0.28046795477615, -0.0592263094975949, -0.133982544951981, 
    -0.25887652048085, 0.281325556634855, -0.226157750761627, 
    0.0455761504543707, -0.0565735020952901, -0.035410574433589, 
    -0.0274329626883704, -0.0228122907871279, 0.0191373551018356, 
    -0.0824492733992229, 0.0322065060606327, -0.0153294321968896, 
    -0.1007165438052, 0.0526681922953064, 0.2135021209707, 
    0.0387073327842285, 0.278259797962841, 0.050122386274276, 
    0.269619829214934, 0.875960622730416, 0.235423895574999, 
    -0.170769448136413, 0.37245855154723, 0.781776635901514, 
    -0.0608873976516047, 0.400564752890298, 0.742627360076667, 
    0.423848840431961, 0.114166429251326, -0.245882066173994, 
    -0.426604760694145, 1.10808707999176, 0.359983074031636, 
    -0.140221528186428, 0.335851830849541, 0.460185211018369, 
    0.37254910017559, 0.201275028530718, -0.293680185926854, 
    0.223490021202593, 0.487710518143766, 0.201779044185997, 
    0.0765283957148935, 0.0773640103586576, -0.0252637403393108, 
    -0.17832009889763, -0.273990797557309, -0.0561051485556752, 
    0.0301001800562802, -0.0959558936701967, -0.105918349805861, 
    0.27989492915903, -0.0809511781083954, 0.0792956710869479, 
    -0.0610012116076117, 0.0914608847384713, -0.0627227689795827, 
    0.05161094302865, 0.0532657730090051, 0.0952358644756241, 
    0.0451026308581223, -0.023942617716294, 0.0561338817933882, 
    -0.0184983875503485, 0.0315343282972957, -0.264304601687064, 
    -0.00913633638431158, -0.0941329928314009, -0.20180224587697, 
    0.13571605526141, -0.06027393304336, 0.105914658129468, 
    -0.166122513800771, 0.0282468354909273, -0.00679777341347465, 
    0.00960591847095498, 0.0373222205279345, 0.0308002069237555, 
    0.0235609743029394, 0.00153381345928826, 0.0933348763842697, 
    -0.0399426941727036, -0.0807827953173604, 0.0981519793805008, 
    -0.052138928611505, -0.087764689273625, 0.666538885280016, 
    0.22790239826096, 0.140534140446245, -0.260325046853404, 
    0.626396479330387, 0.215969591520817, -0.153733400587662, 
    -0.0967883445401283, 0.585256860044092, 0.594379181329616, 
    0.378122317021654, 0.224090363847367, 0.196711383160188, 
    -0.468561025381728, 0.525214278906193, 0.473835593511436, 
    0.181056862325681, 0.046288164605038, 0.331392648962443, 
    0.148766606846175, 0.0734878137965056, 0.0512517725632217, 
    0.08570724965614, -0.08722422957853, -0.0286247745631792, 
    0.311974674330795, 0.279741210269684,
  0.184683846625497, 0.018076986055987, -0.343525238853372, 
    0.416253648487155, 0.476137505965257, 0.258847990201698, 
    0.178528982196878, -0.384824204418659, 0.288042170198186, 
    0.506873496489746, 0.0775818196681145, 0.0890365837837839, 
    -0.192986249395095, 0.300642398606735, 0.251044448137058, 
    0.059870663638713, -0.14485187808436, -0.0275339541249313, 
    0.268291805330491, 0.19016533429239, 0.0355178753225216, 
    -0.0779285171345521, -0.123425104157095, 0.160721846552531, 
    0.277096902030114, 0.0792535806937224, -0.148644035133091, 
    0.0896713686937074, 0.456895466553431, -0.0730156248619211, 
    -0.0685102312957103, -0.0192977640103831, -0.0202777978415258, 
    -0.0293090554788218, -0.00902059338474827, -0.0359173688785552, 
    -0.017007392429807, -0.0268032906896476, -0.0104997225923253, 
    -0.0555376253534556, 0.0457039853672508, 0.0709408224942137, 
    0.0911171856323363, 0.0812716260812374, 0.0863749034016723, 
    0.0723390441082009, 0.0787394485993417, 0.0856212830263136, 
    0.0850274346817199, 0.0502468460780832, 0.0826629338576198, 
    0.118157069516299, 0.171616451713788, 0.130183420018273, 
    0.0593878636898098, 0.248562058818881, 0.194165688116603, 
    -0.0873021292475447, 0.230158420245997, 0.318441069663987, 
    -0.101336905400598, 0.561540029577295, 0.572780454210473, 
    -0.281811701430047, 0.262112953890074, -0.518986797839072, 
    0.906789426386861, 0.176698220579041, -0.236065448848967, 
    0.26795088742035, 0.554750216267728, 0.202831265649594, 
    0.189190261432549, 0.286990296445548, -0.0627473105463117, 
    7.47961561954752e-05, -0.281760133802688, 0.124652481951694, 
    0.00608245490212948, -0.169068016368099, -0.152678658184046, 
    -0.12957029841143, -0.175964228310647, -0.121612736443755, 
    -0.143180519462486, -0.114534401056387, -0.123894487498554, 
    -0.0747251550693259, -0.117011156457041, -0.0207442421263312, 
    -0.100102069318816, -0.0570234306860424, 0.137145437311697, 
    0.396873881499378, 0.303669708698305, 0.115491018978976, 
    0.118074653864946, -0.0997432914768841, 0.599609142050594, 
    0.0416308664885469, -0.0544036683497619, 0.011210820964442, 
    0.454016536236328, 0.212633182797784, 0.425764988789359, 
    0.492661186697461, 0.23844531377936, 1.06360302180148, 0.430137498877289, 
    -0.0469772250796832, -0.160522178508289, 0.0366652153517136, 
    -0.15940197963692, -0.023586438741613, -0.105856910765661, 
    -0.126300527782448, -0.0536825990005478, -0.0872862191941575, 
    -0.0564910527169044, -0.142601883997763, 0.0291371014077759, 
    0.121977804350565, 0.0946504151976062, 0.0684367307469152, 
    0.0646986089627396, 0.0482445377589481, 0.0790478864374596, 
    0.0840818770345004, 0.0511377698147431, 0.0709561084327344, 
    0.0268855830235748, -0.0164296715002717, 0.0630664737627427, 
    0.0176478008019902, 0.041527468458305, -0.0196053413293668, 
    0.0325252360727215, 0.00599582798484383, 0.0474342214208223, 
    -0.0412127338778001, 0.0428354724359666, 0.0869462775559989, 
    0.0814020423858024, 0.13452794284605, 0.171043332445007, 
    0.0768297217391236, 0.0939629924506667, 0.359140829365894, 
    0.044721009602672, -0.248431498274391, 0.0687535479669, 
    0.481079736325129, 0.0828885403017021, -0.318094575212837, 
    0.218428941724837, 0.54312176187989, 0.351329068332967, 
    0.163246362449998, 0.0300051531680416, 0.192262241661075, 
    -0.123070191517538, 0.0461686649512269, 0.409279776320137, 
    0.72591632864876, 0.35665446520356, -0.115506044512285, 
    0.497290563584049, 0.39017008240329, 0.0386778029543979, 
    0.0417545059989292, -0.055689022892608, -0.225488141161777, 
    0.119745513176657, -0.179803064226097, 0.0761426773817726, 
    -0.315760768508835, -0.00948179669485783, -0.197847344628815, 
    -0.014618649687653, -0.339794129498485, -0.0784405993960755, 
    0.0711833221522492, 0.155973478868775, 0.1257223440515, 
    0.112680455478364, 0.107711330853905, 0.129724525903466, 
    0.167964962737786, 0.14711504256155, 0.0928808855953361, 
    0.134064457741777, 0.13693023413146, 0.132953237305013, 
    0.200114480170766, 0.255014624408156, 0.191761610302464, 
    0.134081251337102, 0.260102651910711, 0.335001614256449, 
    0.199527116502858, 0.0677005410899547, 0.0611010816351655, 
    0.464776555356794, 0.381968420033252, 0.112712032411452, 
    -0.143453142877367, 0.11987173867659, 0.34524103741478, 
    0.367448819035343, 0.622541576237786, 0.26477463553816, 
    -0.321526761374623, 0.233314344444747, 0.518021898881879, 
    -0.0350318773411234, -0.00169843299795637, 0.0174372215937534, 
    -0.287974934369489, 0.225819865007057, 0.569454604393216, 
    0.285479100249867, 0.129632991970979, -0.114500579334576, 
    0.329792071663492, 0.160455854161788, -0.338023828680867, 
    0.396583528465495, 0.181035801047018, -0.2513337347511, 
    -0.16275563000272, -0.257599145732999, -0.230829032668523, 
    0.0273522596472135, -0.0660613908636404, 0.0918797273236923, 
    -0.273247775764775, -0.0400516206307585, -0.102275867223335, 
    0.0128325429590326, -0.285145814003304, -0.0140243690561337, 
    0.0843528571317492, 0.0894196128756241, 0.156285367383848, 
    0.191098876726108, 0.175216017907017, 0.214062201874674, 
    0.24844850932352, 0.15698951888301, 0.0209723931470456, 
    0.0492205559242982, 0.489749332020974, 0.316114296151104, 
    -0.0156141415335983, 0.181125974254923, 0.627001949677576, 
    0.274955169403705, 0.0590426895960493, 0.359093605046964, 
    0.314825525354125, 0.27241541861611, 0.660453835344331, 
    0.397376285719074, -0.0677181545225375, 1.12890354552824, 
    0.51494402260422, 0.0271857206492703, -0.216644092821006, 
    0.23330810454362, 0.408095111017376, -0.206400937320844, 
    -0.0426779428729705, -0.117760851807042, -0.0849058115031108, 
    -0.113104132274899, -0.102769137494214, -0.0904905651254441, 
    -0.10661832109093, -0.0533064003709473, -0.118871029477091, 
    0.0477209168178801, 0.106662364513129, 0.122779175538973, 
    0.123224121207144, 0.130656698032726, 0.137520191241355, 
    0.139244187429369, 0.120059583773158, 0.133971219877068, 
    0.14498779497697, 0.11596360857515, 0.118035686481152, 0.114119969632897, 
    0.110468338157651, 0.0763027305633191, 0.0723337914462383, 
    0.0907015777846715, 0.128327674670392, 0.121696530484948, 
    0.00774439923575144, 0.108451150642943, 0.150625493631924, 
    0.305083141442627, 0.412027567403236, 0.147447858624605, 
    -0.12508644074127, -6.74280730011551e-05, 0.536611286051499, 
    0.310209570828477, 0.230584787447303, -0.183497118264284, 
    0.680673674047112, 0.173637569427904, -0.314092579259275, 
    0.00717710742809953, -0.766239572019292, 0.862678639888302, 
    0.260912814432249, -0.0942883080215628, 0.369047374734837, 
    0.396415489656591, 0.049523768194875, -0.0146842221090559, 
    0.290750929417445, -0.0321372171317205, -0.0804740703816712, 
    -0.528172769554089, -0.339799560487498, 0.289769882103278, 
    0.120257556502331, -0.0297802357425841, -0.001333879240042, 
    -0.503775298800364, -0.00293762625064337, -0.392124876419227, 
    -0.372411489149731, 0.241576920368923, -0.381655084848161, 
    0.11335698793888, -0.34965177518324, -0.125537985303756, 
    0.0425494263347398, -0.0224333817347706, 0.0138311473316549, 
    0.0184758506169517, 0.0729461618580545, -0.059473191652614, 
    0.0508836653008109, 0.0150539911319907, -0.0369779028425494, 
    0.128757203205656, -0.182191766634413, 0.2354217900989, 
    0.413933333432815, 0.173129549761647, 0.0952483012646458, 
    -0.194208950945328, 0.153704244395814, 0.369453090929895, 
    0.391705572250613,
  0.0781415885602084, 0.0921377271023371, 0.131826056767396, 
    0.22968832713915, 0.200300102879196, 0.0766663920069795, 
    0.0982195482635085, 0.433654810830234, 0.0456157940125603, 
    -0.153785735216091, -0.241840353229945, 0.533194469056102, 
    0.43191421721398, 0.135959128437201, -0.0467323242684552, 
    -0.128149633641182, 0.507799794897138, 0.0277521384954819, 
    0.145358445959038, 0.925850245148217, 0.257096179491205, 
    0.0383853982113913, -0.0345897776471442, -0.105470773047693, 
    -0.0909243400004271, -0.0342484769211568, 0.344710225219127, 
    -0.0528038733969377, -0.0763960738760009, -0.0102250815008135, 
    0.0608443573527939, -0.192776619211845, 0.165491526946456, 
    -0.158248644464713, 0.0892711971323122, -0.164008291247291, 
    0.0756872533161156, -0.111962568311132, 0.110923539373321, 
    -0.302529898323629, 0.0164124742874463, 0.0971640533836602, 
    0.104458708052872, 0.0983898126820206, 0.108398750623064, 
    0.0987045848928581, 0.121377652168587, 0.141185502894376, 
    0.101522253197348, 0.0408714345278733, 0.0837341865255122, 
    0.102777551115792, 0.108728156626733, 0.110995006144007, 
    0.122305225224671, 0.181068584655049, 0.132138344837858, 
    0.0175062217723311, -0.0955390890934378, 0.295120159407766, 
    0.340779797737089, -0.000343803401480103, -0.295701074756159, 
    -0.13517672372929, 0.822965442536472, 0.232838367804305, 
    0.154327472130598, 0.209123424086433, -0.29602485710113, 
    0.00778595908189917, 0.781976176912936, -0.0229168204331632, 
    -0.118305586098988, 0.029295651938668, 0.109308752363917, 
    -0.0100452408144144, 0.745558606160276, 0.575733625915473, 
    0.350877424136234, 0.518044295328498, 0.19428083692478, 
    -0.0507565219688214, -0.0472016694648689, -0.0407782696515741, 
    -0.0415772165439502, -0.050858495214566, -0.0679220969912106, 
    -0.00611048687780055, -0.0850965633141881, 0.059850121001535, 
    0.335109051484335, 0.000423955867255535, 0.137598221282583, 
    0.272974205864302, 0.267657567321797, 0.543236447345501, 
    0.340469345126046, -0.0913498961633079, 0.512263911884411, 
    0.44454206002049, 0.00622414967741199, 0.17132479376161, 
    0.700031894626219, 0.313388194262389, 0.185323820661156, 
    -0.277532731819813, 0.0844872470420567, 0.480223213761666, 
    0.359268804667342, 0.245504279494556, 0.141614424410695, 
    0.0733020465830909, 0.289139274020854, 0.486849010693879, 
    0.212207486092539, -0.024623377397784, 0.191058711091628, 
    0.407815813791402, 0.190159532448868, 0.164210334834823, 
    -0.253378666330812, 0.112996162705311, 0.402756632289209, 
    0.398854117162565, 0.261454143184274, -0.163920154392988, 
    0.420655218339836, 0.457231670314646, 0.267655486514542, 
    0.163739806014542, -0.234873764365304, 0.382809757853345, 
    0.274082650407232, 0.102285547895297, -0.220105781469962, 
    0.423027472093485, 0.165326568195695, -0.105504883778059, 
    -0.0116840750866058, -0.0335795029419619, 0.0955229987072389, 
    -0.125850054550873, 0.117562491846851, -0.101405538094462, 
    0.113097493836609, -0.102852784813848, 0.0851045331757877, 
    -0.196060730309974, 0.00574148076296488, -0.218694387563795, 
    -0.0934496181225664, 0.0622865159487598, 0.28742856004129, 
    0.143927101004013, -0.0237569751018228, 0.355955546854938, 
    0.43813222814128, 0.181640385628851, 0.0431972438336128, 
    -0.000160687932402807, 0.316675187727954, 0.492527523288087, 
    0.377107550550902, 0.30373924401032, 0.346164579484651, 0.31733707274206, 
    0.270134620551087, 0.341920847460826, 0.317407584857613, 
    0.23028716108951, 0.362668346238341, 0.39465279912267, 0.152983499440334, 
    -0.0897566034296631, 0.351901256526757, 0.444657689250259, 
    0.153001442622256, 0.0697547635677416, 0.194101564005261, 
    -0.010551223348369, 0.749492628296746, 0.0753025043105817, 
    -0.080502560247907, -0.190591307728025, 0.564316253967401, 
    0.33354158224059, 0.118741687732923, -0.270800047238775, 
    0.22822120999911, 0.406351375383104, -0.31954540530872, 
    -0.120707379875258, -0.158108804695434, -0.101420894169283, 
    0.0362295058085739, -0.161042042808465, 0.0450158643377289, 
    -0.0147873894737776, -0.0223322804500622, -0.0313161343635892, 
    -0.225244641878921, -0.0711273486348714, -0.0499120608245673, 
    -0.0622589464941819, -0.242436974937443, -0.103316434774863, 
    -0.0905339142490574, -0.286473540575666, 0.197401567869927, 
    -0.08256360308328, 0.145771125040145, -0.0252854254427183, 
    0.0243609035141782, 0.00162024225233459, 0.0319415750783083, 
    0.00567379788510937, 0.0345554046114939, 0.0170736691053803, 
    0.0232307678629346, -0.0790639957956017, 0.0156130683395648, 
    -0.0109915155656739, -0.00439384396282541, -0.00211930497997458, 
    0.00321043833919619, -0.00721140523595057, -0.00798565542023563, 
    0.0899144371369728, -0.00078258139377102, -0.0372870906383181, 
    -0.202205020326015, 0.463039572601581, 0.201226014095444, 
    -0.135673820577568, 0.496669625259359, 0.432593588692023, 
    0.188820183437719, 0.379972743741049, 0.395145688793279, 
    -0.430533270636952, 0.162901844649545, 0.863269989655849, 
    0.290285204135594, -0.274171402471218, 0.424536506768335, 
    0.628223715059197, 0.325038295544615, 0.150656725057342, 
    -0.137056421949549, 0.188924315990195, 0.681593943074261, 
    0.0792146771173392, -0.0964607618356671, -0.0539779311521853, 
    -0.0581586348117506, 0.133829878592636, 0.031789945897535, 
    0.0186532762688659, 0.0564775362141452, -0.184105608052979, 
    0.0456275868062605, 0.1696731928535, 0.218549562488572, 
    0.144238606957996, -0.0299886895583451, 0.16256684919788, 
    0.214010842282834, 0.102275116233235, 0.139533330591833, 
    0.253055632461097, 0.0409791574937162, 0.0084762359181324, 
    0.0132020772869914, 0.0482065614817865, 0.0260652097908308, 
    0.00195211445972886, 0.0287975562709948, 0.0320471677736155, 
    -0.0463155914799397, -0.0304070689517455, 0.0127863739261943, 
    -0.098565490885235, 0.047156519490612, -0.0686087948294, 
    0.0297060015722229, -0.102582000795125, 0.0145559148487697, 
    -0.0599851515091547, 0.0189027229374182, -0.123445354480971, 
    -0.00325448343144483, 0.0473831539146633, 0.080885530494269, 
    0.0831403265794667, 0.0799295019970573, 0.0856532646930399, 
    0.0972912138856247, 0.119363099949585, 0.0905813198266987, 
    -0.0529541694132096, 0.219409064269645, 0.198075345920677, 
    0.100666002763872, 0.488003473780615, 0.305288978650861, 
    0.0493851321486322, -0.0833630930644251, 0.500353329901521, 
    0.308937441316315, 0.43942526561132, 0.343296947879243, 
    -0.00135153683724235, -0.477228264739606, 0.717745193799907, 
    0.3876384385847, -0.00527519694055804, 0.00746176863284373, 
    1.13354397245914, 0.206073139701794, 0.0607141808162125, 
    -0.272683228590109, 0.0989629837798638, -0.26187336699877, 
    -0.0904076844837804, -0.17566205319622, -0.119606331105239, 
    -0.263740324630132, -0.0934686724709789, -0.26492910192033, 
    -0.0519167629465955, -0.104279139037982, -0.0957688802028672, 
    0.0841411843838002, -0.0694444571142509, 0.0814916579231658, 
    0.0340416567902746, 0.103541214183369, -0.083607558062159, 
    0.046988124608812, -0.0663896066259966, -0.0525786870473856, 
    0.135980203962082, 0.19373898018105, 0.0281155717101436, 
    0.341653209908349, 0.341538749886369, 0.0870240640499547, 
    -0.0876020075684947, 0.350110844955216, 0.339381710464947, 
    0.160420639905618, 0.118780350578902, 0.0944734961135154, 
    0.10529231484669, 0.146457896884847, 0.122294076590136, 
    0.0682460086928026, 0.115219769653814, 0.090643064604733, 
    0.0638535185853148,
  0.0985477839922649, 0.123221268990587, 0.133371440576746, 
    0.143004290488769, 0.140174750625082, 0.148742905555685, 
    0.185098669697536, 0.143480755281379, 0.0368722882713149, 
    0.0684943841577152, 0.384301831826853, 0.187727305272394, 
    0.0333799047905436, -0.0763666159037786, 0.182398180687562, 
    0.371616133465237, 0.547809079421104, 0.237768939071119, 
    -0.208212795674592, 0.167594501398736, 0.281767911734569, 
    0.253760710586279, 0.602146249950173, 0.326227268605328, 
    0.191934794234278, 0.278828404549703, 0.0552507441801357, 
    0.54375116349677, 0.217135348259668, -0.0366245841040738, 
    -0.140012891363718, -0.270398578671832, 0.12342312576011, 
    -0.0780664471725911, 0.117101177620812, -0.178989588708917, 
    0.0433514977114164, -0.121051975635666, 0.0261790979249949, 
    -0.256559132185976, -0.0283499313245114, 0.0688655285578475, 
    0.147944465494499, 0.165730715152741, 0.170847656932973, 
    0.140205204618628, 0.122558465337441, 0.162747958464949, 
    0.181851369798525, 0.142148021602365, 0.147974352314114, 
    0.153890608629324, 0.158768538528198, 0.192989159102897, 
    0.204906720650458, 0.16465627275643, 0.175025746616078, 0.24703261905962, 
    0.189915496236302, 0.121802725041703, 0.191034312382567, 
    0.148543198264093, 0.314782500613077, 0.400895792241765, 
    0.119151226661048, 0.0431155327793673, 0.651769265005031, 
    0.381296788626991, 0.0988795871859595, -0.196473406281537, 
    0.0806984171054252, 0.257924425713029, 0.352356487584883, 
    0.669442815764955, 0.265409555767614, -0.4201346628131, 0.19602201864135, 
    0.885142780892988, 0.0141803238436049, 0.043550019830226, 
    -0.196361388866124, 0.00111312737856559, -0.183703608891067, 
    -0.0567976983510329, -0.0183276598678375, -0.0544140027933497, 
    -0.000690717266499552, -0.0758777074070424, -0.182321379793962, 
    -0.0155013844815874, -0.205881269166992, -0.118457973288243, 
    0.0316881913135114, -0.0363104550678412, 0.122844754373232, 
    -0.205986965728637, -0.0168759541734781, -0.0573146356591899, 
    0.0642926423839584, -0.0632408913913728, 0.118704578652731, 
    0.0119301992380629, 0.0845464273493037, 0.151834829519957, 
    0.0653678398277013, 0.107240015288191, 0.12911316699367, 
    -0.0420939551239539, 0.057128400734697, 0.375972985156863, 
    0.587106593907777, -0.11540351407118, 0.784660686273028, 
    0.523526446268411, -0.330588831715204, 0.437406191026075, 
    0.813134627148446, -0.075053398503896, -0.0602563428146826, 
    0.0588403573622044, 0.433634372340662, 0.216642940567254, 
    0.0207151951937609, -0.00982639540026327, -0.123544248639151, 
    0.401154324270744, -0.0436098241653849, 0.362250908808055, 
    0.390091956684307, -0.19680034603132, -0.142646054901599, 
    -0.129179341929515, -0.0785402739674356, -0.168268667112994, 
    -0.0229706052362963, -0.100388533257808, -0.0517075269249643, 
    -0.11024620196159, 0.0130665497213445, -0.111779998596384, 
    0.0694469466566941, 0.119427941688713, 0.0922225637101377, 
    0.0435589956801545, 0.143395697428658, 0.180235933372825, 
    0.116036580490348, 0.068811790309861, 0.146473655068269, 
    0.184023614519748, 0.0544010482944429, 0.0704051888535865, 
    0.044717923430391, 0.0479879696653956, -0.095766090990702, 
    0.0116808197489197, -0.00183645953590844, -0.0277284085350124, 
    0.0787633605127525, -0.0501856402538519, 0.042698830250372, 
    0.0814606831859337, 0.0848803101130116, 0.121940402168669, 
    0.131846486191836, 0.0969626682465461, 0.166541773744705, 
    0.207832011043099, 0.118842176830638, 0.10454441053439, 
    -0.194188313217201, 0.214812946052254, 0.245874372006473, 
    0.302238367784943, 0.788009999562649, 0.300374906826557, 
    0.023696614171239, 0.222083984788793, -0.581023170850672, 
    0.356676523566298, 0.523592186994143, -0.0377860672736411, 
    -0.109078478276112, -0.0381861773553705, 0.111344907477231, 
    0.331079636804362, 0.394583361492804, -0.0702823130448615, 
    0.443495458738759, 0.850288890975498, 0.113352909193045, 
    -0.0067906196169059, -0.0103918145201424, -0.00770204296061337, 
    -0.0152512693549706, -0.000559071628120744, -0.056584354392221, 
    0.0533202721038746, 0.186771877781857, -0.16033183592622, 
    0.0470533838937033, 0.409080496208144, 0.216344665682378, 
    0.0787388350240543, 0.532444650064894, 0.308738139093487, 
    0.12776886232529, 0.0999742673267429, -0.165989626971216, 
    0.51621146006363, 0.481964042813691, -0.0551774038512215, 
    -0.207351639811245, -0.0582937174472515, 0.491385349420114, 
    8.04751612568794e-05, 0.29883287211406, 0.836402560592505, 
    0.506965783838753, 0.370696538656489, 0.501049107889164, 
    0.476796977098877, 0.321915152700924, 0.145029758401144, 
    -0.0463457345841662, 0.318906925107833, 0.0369435830483197, 
    -0.0376636878759975, -0.00561427358514546, 0.272842779236999, 
    -0.0764319903396055, -0.0379808156420496, -0.126332655164097, 
    0.0497579525811665, -0.103881424691763, 0.0401969303266899, 
    -0.0176075469002046, -0.192165623119526, 0.0460076067104098, 
    -0.0869930590351771, 0.0886171206946508, -0.118268150323735, 
    0.0717092332961327, -0.0921775406963627, 0.0317662553600744, 
    -0.126166418817318, 0.0369649410529553, -0.100134549667869, 
    0.0767960001351021, -0.183238516193389, 0.0764268328332747, 
    -0.0164368935458793, 0.00942932036588887, 0.255245518164201, 
    0.151742735202891, 0.0489108864524541, 0.32233482198475, 
    0.0192675099818418, 0.0648615696230882, -0.361677328854811, 
    0.462799512447845, 0.330955256472172, 0.0260823940728615, 
    0.785198328372901, 0.492246917427552, -0.190176683165658, 
    0.0442059120333478, 0.704252010078676, 0.345056124213179, 
    0.112255345171861, -0.117550566681292, -0.278255934658908, 
    0.455711194835256, 0.232077420440489, -0.142093687915804, 
    0.455175351729332, 0.359016836663885, 0.0892446502338506, 
    0.481147524761043, 0.293702958811247, -0.165640289191704, 
    -0.0924280175066035, 0.0151218076152418, -0.185150797507617, 
    -0.131599057756711, -0.0867763488385209, -0.0204804542611572, 
    -0.136997176544606, -0.0560932722373174, 0.00802835114054147, 
    -0.0817678544260003, -0.00834819819527329, -0.0134317200343209, 
    -0.0183758001933131, 0.000853007594350738, -0.0494252063642981, 
    -0.0181278444936667, -0.0384682554092133, -0.0401643570379787, 
    -0.0228142313987579, 0.0251249140810136, 0.0170828586909699, 
    0.0363726358331168, 0.0419366558565739, 0.0547167029989461, 
    0.0340068287854848, 0.050996057447139, 0.025041514391379, 
    0.0211667466471054, -0.00152585096448366, 0.230217460058444, 
    0.161536902818206, 0.0549654435518429, -0.0123869723312286, 
    0.447085466324113, 0.364587125559861, 0.170545430140416, 
    -0.102128967210837, 0.720319091373232, 0.178749438621744, 
    -0.160378439187008, 0.528245742895054, 0.379299152936581, 
    -0.105933571077248, -0.393907041120847, -0.0912812288523208, 
    0.702282739645344, 0.941817233326961, 0.0186151494963707, 
    -0.342756127501699, -0.232511180710564, -0.144185951066462, 
    -0.0734999707802787, 0.00520347754258972, -0.0629361949848477, 
    -0.088120378489426, 0.023036241862187, -0.102307887558531, 
    0.0243704225408128, -0.0023868839419377, -0.00220855588022702, 
    0.00991601867490334, 0.0212222093694996, 0.00804230084720825, 
    0.0352333087232078, 0.0249602533808917, -0.000262321842881621, 
    -0.00517117349611013, 0.0508134338741896, -0.00343538336584925, 
    0.031630506711256, 0.0651033991039995, 0.0676151072105311, 
    0.0669145216621012, 0.073336733600824, 0.0639301855569006, 
    0.0682083918773372, 0.0752378821493038, 0.0766077299576939, 
    0.0435464474068814,
  -0.131289864584054, -0.0565555028983443, -0.0836459725598909, 
    0.0507879879376418, -0.0342032253380897, 0.042421880148189, 
    -0.0641664669006509, 0.00864238472201859, -0.165425436003801, 
    0.0479556326332106, -0.111122025398175, -0.109699469516571, 
    -0.257058598137919, -0.133650466597633, 0.00376785162496931, 
    -0.284890538639388, 0.187654574579151, -0.086715499708018, 
    0.0786031665375665, -0.0696971433023407, 0.108279294037042, 
    -0.0318197410895133, 0.0126851427133536, -0.00684563257942214, 
    -0.00647269948579451, -0.000690326333880331, 0.0396321818244519, 
    0.0527098642876693, 0.0141519646533731, -0.0508328628936006, 
    0.0163731699757435, 0.0043272492324659, 0.0232133405874129, 
    -0.00654602674981289, 0.015211232602736, 0.112560217988127, 
    -0.142951611869622, 0.241100372646471, 0.10832710709983, 
    -0.146597372629493, -0.14784151551293, 0.721804620558377, 
    0.0106857727602735, -0.0374545211986456, -0.055032175685416, 
    1.00689199833425, -0.124174889767657, -0.233009329068769, 
    0.513860365161588, -0.066192927260728, -0.179910991531308, 
    -0.536124871552654, 0.280803920804267, -0.0512972910207619, 
    -0.174434504359757, -0.00520554829583289, 0.191792764857938, 
    0.0375114788292169, 0.337271174031985, -0.160373669902302, 
    -0.372623255629957, -0.115551289314289, -0.553769249957311, 
    -0.259259350298597, 0.0496589139519887, -0.598349030913336, 
    -0.00730256870823647, -0.0423277633061033, 0.0936807771066963, 
    -0.334916511059542, 0.0668625916094871, 0.0619657757649325, 
    0.0648038693306141, 0.0949425444214317, 0.103777342434827, 
    0.0686286136427813, 0.0848578921232937, 0.039383990295446, 
    -0.0316990770890879, 0.0711700475427, 0.211686275754365, 
    0.0979914784408251, 0.25062631051196, 0.241021009854844, 
    0.0381693339375255, 0.334133023576223, 0.421535958270667, 
    0.203077022342841, 0.446298605377118, 0.267524062278956, 
    -0.379811056310162, -0.00837641966656993, 0.079073790568885, 
    0.501858826780084, 0.954422193190377, 0.52147047525863, 
    0.665951887230317, 0.801462375642637, 0.357518090270234, 
    0.562349420789256, 0.341796359470469, 0.0578801557050266, 
    0.0071493378154944, 0.0348012881174105, -0.0900940929825924, 
    -0.0216844688398984, 0.162026585628577, 0.0506646953020122, 
    0.176001291687353, 0.247422728877859, 0.0144592068506008, 
    -0.0195060934272859, 0.0538289040495691, 0.0814324758566502, 
    0.0199605375305917, -0.0268446967584742, 0.0418191013263063, 
    0.0660452780596249, -0.0191265753432566, -0.0344198640842717, 
    0.338429478741283, 0.0740868247322766, 0.119416751271709, 
    0.545954453199195, 0.252399194330061, 0.0982806379299055, 
    -0.208781858493939, 0.105522321699211, 0.428332619855837, 
    0.291563876929091, 0.202866949788122, 0.0705930514012189, 
    -0.0989258711278189, -0.225272771936122, 0.529089368529652, 
    0.371228509910921, 0.0809027438575406, -0.068465622104988, 
    -0.110062616964175, 0.280678964915738, 0.330913348279296, 
    0.257361708336762, 0.0653257186568674, -0.0413124441491659, 
    -0.065785215986533, -0.0449202631319791, -0.0554286238092276, 
    0.0562769471714778, -0.173236079917622, -0.154588385188894, 
    0.0387110013118166, -0.11576827609599, 0.0952025348504355, 
    -0.100529176521921, 0.0669024976560455, -0.103961564452464, 
    0.0570536843276098, -0.1429902618286, 0.0237520988995627, 
    -0.111335421258016, 0.00249549872081303, 0.0290574430529275, 
    0.0206676631659318, 0.03495361198791, -0.002696391494958, 
    0.0315842759697177, 0.00977999707140831, 0.0135943468689283, 
    0.0853944538847383, -0.0142420540340259, 0.113722250870675, 
    0.145307783038841, 0.0592769887464335, 0.108693196094929, 
    0.299098116624535, 0.188605128253438, 0.0509517455433543, 
    -0.00615454429630168, 0.356152927354327, 0.257413739324165, 
    0.132794400644599, -0.208274998592161, -0.0101711059979577, 
    0.604100703413943, 0.240618785408991, 0.0466633336021722, 
    -0.204773233658923, -0.0162537997655822, 0.552926992425824, 
    0.408773910585672, 0.187188697917891, -0.194122155780221, 
    0.462430679542048, 0.136450123916433, -0.084917406969126, 
    0.114513262398045, 0.170093630113975, 0.30911104991418, 
    0.537000751427109, -0.0224768623185121, -0.233542329234975, 
    -0.126842274368675, -0.0959871023415612, -0.185747586081691, 
    -0.0851281114647622, -0.195981588496569, 0.0165190787216299, 
    -0.25068888632319, 0.0383321916899777, -0.127064953194614, 
    0.10203668930935, -0.100866573001927, 0.0435587910831745, 
    -0.0286838071592755, 0.0584515810816425, -0.160461971553752, 
    0.0334114588610023, -0.0353983348136014, 0.0449652512665682, 
    -0.150670498174092, 0.00278196424956668, 0.0340506403732352, 
    0.0460160418056501, 0.0476354659268483, 0.0458906065418275, 
    0.0280069754785836, 0.0363824623302704, 0.0435005648777285, 
    0.046063504300978, -0.0207997486446927, 0.0932923171463427, 
    0.149689973729174, 0.0937490811793767, 0.151069658062738, 
    0.247354129344875, 0.125894100514562, 0.160753878386933, 
    0.356944996810832, 0.288976202165831, 0.160610892900188, 
    -0.141385721585552, 0.147514535595211, 0.0663606807941738, 
    0.505227110528522, 0.743246487155789, 0.0758241453322396, 
    -0.0637434755377334, -0.151292752468206, 0.597054697431141, 
    0.151136696940595, -0.0700305332166701, -0.273199404053655, 
    -0.163692820729432, 0.142930715647963, 0.319341680320826, 
    0.189648978812092, 0.10134421296721, 0.190081100211287, 
    0.0628984048539797, 0.0589942999404149, 0.103380093510961, 
    -0.0347497863809694, 0.279818809871203, -0.0619032042604953, 
    0.205683179603635, -0.191727601824903, 0.100678210795154, 
    -0.0497438716684378, 0.152395089566349, -0.21778244946876, 
    0.0866622425101088, 0.0528950945201922, 0.0645532419468113, 
    0.0748806479901278, 0.0704690772677197, 0.0286920732380531, 
    0.0607332645011953, 0.0301305530928692, 0.0298241501371941, 
    -0.0303796228407332, 0.226760853629955, 0.146948424579502, 
    0.0246862987772869, 0.337141603065545, 0.304845647872334, 
    0.125553459914737, -0.0393219614271865, 0.482331381750391, 
    0.187625675460114, -0.232091877382541, -0.23260761655509, 
    0.514424929268456, 0.832728120465295, 0.177200669717956, 
    -0.0789781759155379, -0.255091775877675, 0.404964170446764, 
    -0.124728785736496, -0.143323582207667, 0.652253093996169, 
    0.163783008524559, 0.0103528999317747, 0.203410850708007, 
    0.112828142041431, 0.202008492156883, 0.161108241991947, 
    -0.0488163898228937, 0.193071536263246, 0.00504069308654362, 
    -0.154253426372302, -0.0717517903200168, -0.0606904113596168, 
    -0.0603267080151891, -0.0100012509675023, -0.075756159071641, 
    -0.0196361721993129, -0.0733866446699509, 0.0169656881192326, 
    -0.0445673438729457, -0.10935088539871, 0.00214029493080804, 
    0.159342649014293, 0.0829115725876383, 0.0838731868361999, 
    0.320109255653839, 0.209158659272239, 0.0593663052230446, 
    0.0946908234277911, 0.294929702236108, 0.167774524148128, 
    0.0416070178194338, 0.0213053211882458, 0.0867966503448864, 
    0.0526414933324562, 0.0768094171305116, 0.0416230890050789, 
    0.0753539836542586, 0.0559797741989278, 0.0828111863245662, 
    0.0335332876765955, 0.143627799093546, -0.000417612890843494, 
    0.170451296261565, 0.312172506732904, 0.166185861551373, 
    0.0712306330902959, 0.0351417090094399, 0.0237009644631346, 
    0.480599490529206, 0.249772766674426, 0.123343028214596, 
    0.130537467259768, -0.238806677873361, 0.394579169060172, 
    0.416472405668427, 0.545544118854749, 0.398838428477016, 
    -0.265247164148848, 0.401707106004882, 0.53423043601004,
  0.0912169063877895, 0.112613764489479, -0.0798295187802962, 
    0.300219250387692, 0.397519293022627, 0.0490258297467626, 
    -0.0199253221464246, -0.135670534081531, 0.135829111124249, 
    0.325070344679423, 0.261649769994033, 0.114369470589457, 
    -0.0711223843339774, 0.195931755452824, 0.211897849788324, 
    -0.0237376035566114, 0.396828603714755, 0.427765754495649, 
    0.142267235756565, 0.0685956930765048, 0.319904883771334, 
    0.190644920461903, 0.076284635336803, -0.0326896671072048, 
    0.136641949315301, 0.157492446190418, 0.0357132536286419, 
    0.125312477735683, 0.259037001351948, 0.047424856033606, 
    -0.0760925688847797, 0.00455345421194886, -0.266469817773728, 
    -0.0251113554240856, -0.0510441936567534, -0.145532030319057, 
    0.0156172406700349, 0.0255590436443724, 0.0991853036954798, 
    -0.165130785705469, 0.038765291384634, 0.198763812084364, 
    0.103941880673134, -0.0751176125983398, 0.21635064141837, 
    0.306359591299231, 0.106956053730657, -0.0207088694975831, 
    0.332973613801978, 0.336545283006018, 0.229294650086752, 
    -0.327550871845061, 0.3099958301047, 0.822421094004882, 
    0.181430938718782, -0.243385013193057, 0.0290983279125659, 
    0.582458635123103, 0.363295208319938, 0.201188499440989, 
    -0.175633833431207, 0.448175740581667, 0.339901997293962, 
    0.0862246665549038, -0.0974076585053555, -0.184854891606563, 
    0.415535622385715, 0.297673995437069, 0.228339725798386, 
    0.390710442684603, -0.0329442404969312, -0.101131116036374, 
    -0.120639257172173, 0.00972871574297175, -0.218722159533751, 
    -0.0814083155649304, 0.00318124133021067, 0.032885285080068, 
    -0.109544740023263, -0.0643714454721117, 0.0587977246859478, 
    -0.158302548202869, 0.084723358282614, -0.113127791056589, 
    0.0137170359279741, -0.142381781799084, 0.0183884197900696, 
    -0.100558896184372, 0.0511476459517355, -0.243896261252274, 
    0.0108713624382561, 0.0269049631429538, 0.179470381043801, 
    0.239216442750606, 0.112637847333769, -0.0626609330175367, 
    0.164508618215257, 0.445924918240087, 0.221831636548877, 
    0.0530709410600392, 0.100448070390782, 0.31917727531244, 
    0.228508157239484, 0.156113984785081, 0.660078578886543, 
    0.550844208629846, 0.151707984024094, 0.0927210844372961, 
    0.746843983317013, 0.386574162765708, 0.0582696191876829, 
    -0.0982533222320079, 0.549000007929397, 0.450150496147714, 
    0.117496573542479, 0.0203046439341771, -0.179106656662066, 
    0.52745496330307, 0.401280273342393, 0.218344890318669, 
    -0.18431908418594, 0.347379440771453, 0.307770169162737, 
    0.17512617362629, 0.269718724208258, 0.217854472891922, 
    0.0308738144812972, -0.391502610331163, 0.148949772857993, 
    0.543561364585793, 0.156458592038656, -0.040344601200018, 
    -0.199830074995169, -0.140343211185631, -0.131722183625531, 
    -0.128459225123532, -0.133821516071471, -0.0481370148087029, 
    -0.246082396777212, -0.1235496708862, -0.0194665912957631, 
    -0.126511499959073, 0.0661970448162875, 0.000335103033761636, 
    0.0556676165737544, -0.111943208020304, -0.0165770180779858, 
    -0.0598674742868938, -0.0568535244024829, -0.0575031541875262, 
    -0.0815735421641734, 0.116592425096845, 0.005970197031748, 
    0.114785582609577, 0.194359408322112, 0.077126278594635, 
    0.0999025804040455, 0.178839182533921, -0.148126887785772, 
    -0.0872374199724462, -0.461692092583089, 0.575656585326465, 
    0.466591376248547, 0.232307998571958, 0.735991228474702, 
    0.752316742394197, -0.365282234153018, -0.309126473111016, 
    -0.205508611434782, 0.736171500568667, 0.102518645911126, 
    -0.0646719743258964, 0.277784853455813, 0.400947182958036, 
    0.188796008179059, 0.0468213890556916, 0.00423498882006262, 
    -0.15327647061152, 0.091540141713183, 0.257802876306416, 
    0.0177118345078307, -0.0340045235469089, -0.0759609739028585, 
    -0.0564115896980906, -0.107654481573882, -0.0492496536668779, 
    -0.0680319957791703, -0.135604795173945, -0.0788125388553423, 
    -0.0693557273280008, 0.0130219441225017, -0.0356697837197329, 
    0.103980048428692, 0.20185075321792, 0.153524575808946, 
    0.0941239104276865, 0.0822171696851466, 0.141605936931575, 
    0.23248966107421, 0.161725639704651, 0.0522236714139096, 
    0.0359217124469198, 0.0806304700790079, 0.051642627045925, 
    0.0661955342477987, 0.0453914324921072, 0.0603235823891109, 
    0.0653275839716249, 0.0750533565473145, 0.00379148206018158, 
    0.0957721965054283, 0.126845859900536, 0.0631412768918866, 
    0.165992622849263, 0.303222521366906, 0.154264941919564, 
    0.00591699474957784, 0.0244680448664182, 0.417722721127079, 
    0.199839307787103, 0.0888756434999666, -0.00353929024274371, 
    0.211393059653617, 0.00714968638973887, 0.392460299958738, 
    0.819437322030144, 0.0613008490273514, -0.189537984144358, 
    -0.0235571455278529, 0.520997252394476, 0.144843651126894, 
    0.0490707122254451, 0.00968659423159908, 0.253812494534991, 
    -0.0479781290854988, -0.0954802172053312, -0.189122249557476, 
    0.00900340541108749, 0.0230102955604443, -0.21086891018051, 
    -0.11535688414977, -0.328278069434307, -0.105468365193604, 
    -0.0726937774275639, 0.117207841755318, -0.242847115043879, 
    0.161988237359342, -0.263849117976272, -0.00619680079969844, 
    -0.417213864069167, -0.160108532104527, 0.0667821462161667, 
    0.0634490016845694, 0.0377835723928857, 0.119240924855298, 
    0.130850073680272, 0.146461467832595, 0.248678938360302, 
    0.168875836360605, 0.0182330077739438, 0.280031962085154, 
    0.347778677205609, 0.0464793300422911, 0.188701324028655, 
    0.816586539895473, 0.225653379110609, -0.0782157705691776, 
    0.0244827956471186, 0.756218406997219, 0.139560243020515, 
    0.0395506737652808, -0.0982253187667989, -0.0694296075829219, 
    0.330444285586045, 0.925897366343556, 0.316344635718249, 
    -0.0384132522713182, -0.0609718988043913, 0.354421447895722, 
    0.347652200825776, 0.145518751845008, 0.649365117151013, 
    0.830881402126027, 0.118743896579474, -0.233795900491512, 
    0.0982131555839804, 0.104282932143608, 0.284744286496502, 
    1.34496750173463, 0.0755901267279857, -0.274671507117777, 
    -0.204707184962175, -0.0121998286021795, 0.038572500148402, 
    0.0372818679825939, -0.0502349351407453, -0.0951879885732214, 
    -0.275169809022213, 0.0856895221893192, -0.190904096908731, 
    -0.0324530653468756, -0.038600681731633, 0.141607262086198, 
    0.0119440963765188, 0.218597720712318, -0.0483002608181984, 
    0.233442389392789, -0.205103287198801, 0.182211817163296, 
    -0.227312768604879, 0.116947695346213, -0.044678772295278, 
    -0.00997908714881825, 0.251188158600389, 0.143378329931462, 
    0.0308272508926168, -0.0865453378658147, 0.245458163254371, 
    0.269723837570299, 0.0340155886101804, 0.0294488156945441, 
    -0.213400538867414, 0.490636772641403, 0.364984570014373, 
    0.106220465091505, -0.0624730486237375, -0.081534720810031, 
    0.259988407405514, 0.557885877367547, 0.467718906873378, 
    0.18551559379411, -0.0272342289322826, 0.0262795033883278, 
    0.633571734630124, 0.280519524804012, -0.0112069060403574, 
    0.0959480919886437, 0.555118013163729, 0.253317296754619, 
    0.10039269329124, 0.0433134594726913, -0.0840096541979681, 
    -0.0251858312715897, 0.706804296438726, 0.179645893963879, 
    -0.00023116892167438, -0.0934971761326184, 0.61106207843512, 
    0.126530848739038, -0.0503595714736364, -0.117953129609288, 
    0.452189472531349, 0.367940247844595, 0.147626344033789, 
    0.0473983131334001, -0.22496902677029, -0.0829347476991902, 
    0.428667556970999, 0.373524128763217, 0.194447236225912,
  0.103926502399894, -0.0254692205707991, -0.411865775650116, 
    0.579662470959305, 0.451321926983383, 0.111338460612063, 
    -0.0198366292134185, -0.0334978381934809, -0.0690097958134958, 
    0.322451746183326, 0.595743568911102, 0.331129920935332, 
    0.06794768484589, 0.0411518745267059, 0.0899335889029497, 
    -0.205339051049497, 0.073034260528199, 0.293185653897432, 
    -0.0304221007589111, 0.0504097805385984, -0.128045801142884, 
    0.179943718301872, -0.26115651949629, 0.112318700954299, 
    -0.2668902281507, -0.0384910229573375, -0.0797855768468705, 
    0.034689085708022, -0.358254888792079, -0.0659891858688862, 
    -0.0594536057703871, -0.16568485088942, 0.00705830793303755, 
    0.0105812386872106, 0.0354258853413929, -0.0891340820042857, 
    0.0281654232270866, -0.0433026465198122, 0.0224731014437584, 
    -0.270477945721312, -0.00700278050616365, -0.111784752485772, 
    -0.0867179877606101, -0.0626931624873441, -0.0544624741525258, 
    0.107201238649221, -0.211882193905164, 0.120434776625167, 
    0.0695270175610713, -0.325062193971731, 0.0286894113316892, 
    0.345960209049974, 0.0432221915869218, 0.0416697869366744, 
    -0.111712840316551, -0.236238839118141, 0.593673728341498, 
    0.159012700202543, 0.0538293634864358, 0.00181057436263815, 
    0.298259384620019, -0.105711540264649, 0.972471356685081, 
    0.602094440454442, 0.125786368993877, -0.0275931599620719, 
    0.404474825017495, 0.361874977921342, -0.0537638623603209, 
    -0.0903875625522114, 0.483078394032314, 0.320989171636322, 
    0.123994378897845, 0.0795617944878782, 0.0670219729171013, 
    0.0365078516586604, 0.0441636223857961, 0.157219404683246, 
    0.0844782325858922, -0.233969107347647, 0.105285013416337, 
    0.391308666410447, 0.0532255873632633, -0.112999212316231, 
    0.0831046961470621, 0.390643290280184, 0.496132372564329, 
    0.203963601390224, -0.0737500807632748, -0.13766316601192, 
    0.592163270059622, 0.46021178713508, 0.120138977333508, 
    -0.0369824373761534, 0.28973474840182, -0.223922821307466, 
    0.29060724432807, 0.754459685719555, 0.211323992302724, 
    0.0597160486889762, -0.0304866412982965, -0.185532905825698, 
    0.0676865944062303, -0.0507349565903818, 0.0663444104042329, 
    -0.189320332682707, 0.0129863374045635, -0.0311566983394171, 
    0.0976156193769634, -0.192665003267685, 0.204136466105686, 
    -0.0766572119917836, 0.182934922360236, 0.436081326287843, 
    0.177846292220082, 0.0866063798562068, -0.283572886881892, 
    0.0940914791422094, 0.503876589405835, 0.19697915045104, 
    -0.040722987939601, 0.13012573813326, 0.671856361592585, 
    0.430684334581437, 0.0901211821389649, -0.455637038012603, 
    -0.0843995543941274, 0.82845841009009, 0.335930614709463, 
    0.072230165944135, 0.670079861236169, 0.442683564018584, 
    0.0292079590761274, 0.393732806818307, 0.588223205553416, 
    0.260122996143871, 0.189797264954308, -0.203098174173622, 
    0.250820647072392, 0.34533333331712, 0.361333662254821, 
    0.248562622020879, -0.154349838560289, 0.376979010656548, 
    0.260990997626648, 0.0458784124936391, 0.148459236621918, 
    -0.276557904110715, 0.37576262908394, 0.678433894834605, 
    0.0713517415487918, -0.035391276683808, -0.0128290923485135, 
    -0.0532321061662673, 0.0857253148972936, -0.0441823050592264, 
    0.118560535619234, 0.00671166516468484, -0.123405707017958, 
    -0.00536798523575691, -0.220454417241416, -0.0831411639997334, 
    0.0255154634294162, -0.130191693126554, 0.120722593879558, 
    -0.0344130598073884, 0.0921827724207254, -0.060238216960123, 
    0.0656622566567842, -0.165569223076437, -0.00991775716175253, 
    0.0622474756419021, 0.0970193848185543, 0.104296359581852, 
    0.111211305644561, 0.103894264208815, 0.111026221074075, 
    0.137637958343531, 0.118966118991866, 0.0755449854651926, 
    0.148709034099153, 0.170628433467058, 0.172527632370033, 
    0.244829873195182, 0.261140550793671, 0.166068606026335, 
    0.195009771478231, 0.372552646851351, 0.25844579267331, 
    0.153783333937579, 0.185974766688097, -0.294868035970427, 
    0.385839118638872, 0.603158202974188, -0.0573320427158525, 
    -0.160635991193475, -0.0495118007835622, 0.483029830766391, 
    0.165625568185619, 0.374359755660062, 0.246702322813726, 
    -0.321638792328781, 0.18699079723446, 0.364519685390538, 
    -0.271502736360903, 0.0136725705256115, -0.0492212300605095, 
    0.429270729535247, 0.0827360668163854, 0.0860233750870763, 
    0.0190304516938219, -0.255813088877871, 0.189408984298017, 
    -0.16135898223581, 0.038742732366712, -0.335218613858223, 
    -0.0569961563314167, -0.147264964284546, -0.0131591082791966, 
    -0.392372207772867, -0.0674822815688887, 0.131163895220392, 
    0.0980118146929238, 0.166895035083085, 0.285278320706777, 
    0.214741767914969, 0.158442529486651, 0.2591140785553, 0.28762071365879, 
    0.230725755805862, 0.241400086844507, 0.212179516854159, 
    0.223427996818685, 0.350092850716826, 0.283361592011787, 
    0.127008133953769, 0.33698366226592, 0.476015604899687, 
    0.191504583894172, 0.0211163133842614, 0.0199976929036733, 
    0.0913144988144755, 0.596179943660261, 0.527251634815882, 
    0.420086980968847, 0.22659921439649, -0.328809626777428, 
    0.0111566698297626, 0.499286762446701, 0.226794356503079, 
    -0.0018964936503169, 0.184329824848906, 0.271140650769477, 
    0.101756094508422, 0.0207564372233876, -0.0562104148402201, 
    0.155943521743681, 0.184029078379811, 0.10046110941188, 
    0.137301235946313, 0.215830582475624, 0.195233350992415, 
    0.165210371816777, 0.181517446411139, 0.152601479834252, 
    0.0818244103211983, 0.103267108783306, 0.194694201578966, 
    0.0979284023629101, 0.0579648778064817, 0.365258804250804, 
    0.213822992796209, -0.0896365933011033, 0.356281583922532, 
    0.440650388485688, 0.426359993406868, 0.264446732190485, 
    -0.142841507824347, 0.300869581244633, 0.383132240785035, 
    0.239955934082007, 0.275131615182887, 0.232130003627868, 
    0.0418627422980006, 0.734045717746941, 0.0314533397639887, 
    -0.236870932299874, 0.205973054187012, 0.411849346321755, 
    -0.0145093693246053, -0.126547171909261, -0.0109711563813754, 
    -0.151828931099117, -0.103833757442917, 0.0216117295331523, 
    -0.101585244629296, 0.0270201062233388, -0.0470586724089691, 
    0.0410769494062575, -0.131827813607903, 0.0388263109262859, 
    0.060451900152959, 0.156067716360472, 0.288477505917282, 
    0.196683861863932, 0.105955641875293, 0.384432233057976, 
    0.273290790531914, -0.0621935725473082, 0.124963375276679, 
    0.610334767733945, 0.150388090746494, 0.296879189628806, 
    0.932102393457103, 0.252868300868197, 0.0481135274984438, 
    -0.138212617883976, -0.242763092458916, 0.772323262360349, 
    0.174833249772561, -0.131841191138252, 0.0880294457027931, 
    0.373179383467903, 0.127032222705949, 0.0394067202239622, 
    0.0873311190168366, 0.281701575087206, -0.134121144733156, 
    0.349855921726413, 0.415024977075022, -0.0166260919591165, 
    -0.0235543728304827, -0.0997746592879428, -0.177918471072813, 
    -0.187090552649252, 0.0380000752719657, -0.193762250838938, 
    -0.0372966125542629, -0.0591573527984574, -0.114242931205724, 
    0.0303019000022712, -0.117349874465106, 0.0506822549773362, 
    -0.039855781775521, 0.044086925660703, 0.0136520555531443, 
    0.124293387406568, -0.0700778726560475, 0.127516482544579, 
    -0.104674598240427, 0.112173035393318, 0.0602566507685197, 
    -0.0362075434067384, 0.0747956648452488, 0.134617151333797, 
    0.328554607816792, 0.140574918328712, -0.188309875203988, 
    0.0428143300447818, 0.316773889457865,
  0.36703832397485, 0.109346836348464, -0.0792871463102407, 
    0.275690160316909, 0.217852259553593, 0.158698576632039, 
    0.357481005544611, 0.152179225484667, -0.0259199192187783, 
    -0.216186214361882, -0.000965258130046047, 0.497697627195246, 
    0.14265793850067, 0.0240964658664202, 0.140958312546114, 
    -0.180219156382697, 0.279148352116081, 0.500045473209336, 
    0.00650602892991017, -0.0465328801500149, -0.173742932789587, 
    -0.0710073578919566, -0.0381651180252428, -0.151682288863487, 
    0.104284949473542, -0.118906485334967, 0.0109570664910608, 
    -0.0676658186897032, 0.0196067247703966, -0.164742099782592, 
    0.00457733445206871, 0.0794431118737673, 0.0724897870746119, 
    0.121730728356772, 0.202364561616403, 0.132056191394448, 
    0.100837937668886, 0.259853145417774, 0.154340397788259, 
    0.0239097149787546, -0.0846168552058212, 0.556405935158724, 
    0.308222145464009, 0.0518832073882797, -0.116763113172169, 
    -0.227780725812942, 0.634592101458385, 0.286912949511176, 
    -0.129213752041387, 0.431998987288461, 0.469048907614086, 
    -0.114584048466943, -0.495670601687356, 0.00341529207986468, 
    0.676311537160111, 0.210060739642982, 0.0301854240708506, 
    0.0731778334028834, 0.190042205833007, 0.510248599597587, 
    -0.301527951017342, -0.363966242891007, -0.189091968172597, 
    -0.285328326450182, -0.119372598518558, -0.319927738351691, 
    -0.159170467075986, -0.214614446254686, -0.172931471972158, 
    -0.202056919227578, -0.0157107282960443, 0.061365330401817, 
    -0.00270663954375734, 0.0656632091125902, 0.0510599169528207, 
    0.11543919194515, 0.0183688304466241, 0.0661652679801503, 
    -0.0565134706347929, -0.0170424035700135, 0.0348078167907277, 
    -0.00123825378409308, 0.0490774684582099, 0.00950334595911699, 
    0.0334253897333469, -0.0164529365827402, 0.011553140870157, 
    0.0124627679247847, 0.0295808135340472, -0.0410911634348718, 
    -0.0117222404916136, 0.112565662364647, 0.181111140414564, 
    0.110461323350192, 0.018014674712464, 0.166510169025892, 
    0.312970173614906, 0.0913467187740573, -0.0157844797402072, 
    -0.200026228055828, -0.0886439110611743, 0.619345635236814, 
    0.226868933750722, 0.0843596917055999, -0.132835682323506, 
    0.740887778892619, 0.0342481194491032, -0.422046764286866, 
    0.110692193036852, 0.554853712576441, 0.174796385358793, 
    0.194569881260278, -0.198223247037403, 0.261677286665282, 
    0.188613466999553, -0.00149763157367144, 0.251573568197919, 
    0.239131112064718, 0.270381604353116, 0.131496921909199, 
    -0.143622927132644, 0.0756923284871662, -0.46855324268679, 
    -0.0978839069052167, -0.14389927869028, -0.26840381327362, 
    0.0543373697573871, -0.239858206607387, 0.0598864281697503, 
    -0.238338962478185, -0.00532675204422409, 0.0706070101652158, 
    0.0863071658401034, 0.137390192895472, 0.151764673729425, 
    0.106059921686434, 0.109069282384166, 0.189680713201517, 
    0.121506590738234, -0.0421565963436342, 0.0262072804715928, 
    0.405979513774035, 0.305013231630819, 0.105979783212487, 
    -0.0461914660632777, 0.167449619353124, 0.516770058686432, 
    0.365455585063362, 0.130236531433616, -0.279021553798805, 
    0.453753609160446, 0.510182004976439, -0.459559204752817, 
    -0.0127732887958612, -0.255930372754103, 0.405307914477043, 
    0.287439792515559, 0.584983765079483, 0.372796117915028, 
    -0.402739732859151, -0.304942073074947, 0.0257387782153232, 
    -0.17863274237762, -0.149745862752542, -0.0454641567787154, 
    -0.151217514796349, -0.0085766126493429, -0.143563744496638, 
    0.0248273075472296, -0.169417500919206, 0.00376097502958105, 
    0.0910262074488796, 0.141246286594649, 0.16930806004318, 
    0.191753708172676, 0.154147232076322, 0.128680057974667, 
    0.165577080367649, 0.190289081588994, 0.155495785194707, 
    0.156467533992866, 0.160637995274934, 0.169483885246571, 
    0.194906953950447, 0.193749924089896, 0.165355229400145, 
    0.218787188448059, 0.278874836612279, 0.160080010803918, 
    0.0101872422511514, 0.355764141134234, 0.344120864561087, 
    0.11205179060049, -0.109678843487197, 0.301343609323525, 
    0.386807899496622, 0.243480647575768, 0.274172309652102, 
    0.249663138795556, -0.19519260253918, 0.412508533035093, 
    0.46112367481803, 0.392075539790492, 0.313738255107169, 
    -0.135027058683284, 0.397154746717607, 0.531165271177791, 
    0.205469360760719, -0.0963780666053738, 0.22021011545234, 
    0.304185469536842, -0.0215984621829678, -0.132325429892263, 
    0.00731706824522659, 0.164462680332271, 0.0224454483193339, 
    -0.0401615031930937, 0.06498937489394, 0.0547461360498455, 
    -0.0385601846176071, -0.101121953069419, 0.0539763720714263, 
    -0.108402523976153, 0.0144071461491185, -0.182831573165311, 
    -0.0557758925058934, -0.0702224373765346, -0.121307222676525, 
    0.00959905771131481, -0.108065963026592, 0.0508628510219011, 
    0.0959497873140475, 0.125013994834553, -0.0406089970421383, 
    0.36279877635465, 0.25092181280889, 0.00503641059149779, 
    0.065469287336499, 0.483887868575089, 0.0331288473115949, 
    -0.0555720495380875, -0.151264771651788, 0.177446578649543, 
    0.314641310438817, 0.456525016584659, 0.216894382701016, 
    0.915878668981809, 0.924212119910565, -0.00525131647032608, 
    -0.0443094359936265, -0.233216404404623, 0.202512636159328, 
    -0.342809799161648, 0.0855390640974571, -0.444245991730671, 
    -0.110791627694049, -0.287025253140366, -0.169018716130288, 
    -0.217351760980379, -0.132809069865802, -0.0198017093570966, 
    0.172633746103276, -0.0354235326716135, 0.0275487936668766, 
    0.0905644709852099, 0.0838739974753337, -0.0433995981666163, 
    0.0777338317528311, -0.120278254524226, -0.0561473709500225, 
    0.00654749006209539, 0.0880272386645783, 0.0405925976930506, 
    0.0409254733205161, 0.171348692283137, 0.101439663776778, 
    -0.00404242393471031, 0.20201571013466, 0.123311393471338, 
    -0.0802111115667435, -0.333713400422605, 0.508051012396802, 
    0.467098636019624, 0.291361752713401, 0.110770867941376, 
    -0.334509245102281, 0.0140396905602757, 0.689546799283573, 
    0.218055608415616, -0.239960166097524, 0.298089638096998, 
    0.513620511866585, 0.0894100297346591, 0.0664716774012819, 
    -0.336422592946216, 0.671924084142817, 0.299957014533432, 
    -0.119304671677875, 0.384621380015944, 0.453611056981063, 
    0.0365797074066155, 0.0846930419146162, 0.051347980019956, 
    -0.0726131519345151, 0.0631518272179567, -0.145989514183877, 
    -0.0689768859591955, -0.262861752579407, 0.0213906787883745, 
    -0.23933350765227, -0.235545013779726, -0.0738092989330299, 
    -0.0569638878014612, -0.17529942063906, 0.0742228486223478, 
    -0.144935215520364, 0.0825270267519031, -0.131956745116808, 
    0.0737705517346559, -0.119562885607687, 0.0575410647706585, 
    -0.0499616504029123, 0.0221643204310965, -0.0646292900689026, 
    0.0126346641886556, -0.119574683203724, -0.017532491078246, 
    -0.0675304074921502, -0.058718538543079, -0.00233111052863193, 
    -0.0788537263114041, 0.04467548252427, 0.167351043722049, 
    0.248304804382595, 0.116807365942767, -0.159134994786368, 
    0.103842643407289, 0.352614148481339, 0.0240366396562769, 
    0.21310117102321, -0.315915049206532, 0.0711134948526066, 
    0.515216478085146, 0.357094590098939, 0.144253293715917, 
    -0.316100277422971, -0.0157139177197247, 0.532662657582413, 
    0.462663377765562, 0.203619203120618, -0.143245127422945, 
    0.19784597925614, 0.425289676134719, 0.221274958392065, 
    0.144318924558007, -0.174540228250022, 0.323624627308954, 
    0.253518373928368, 0.0257701869017291, 0.281525434516351,
  0.335466155224967, 0.131567069816548, -0.219750706435059, 
    0.025831806905485, 0.430223161165189, -0.000222712027888886, 
    0.600611769890654, 0.745530688721981, 0.137800246224418, 
    -0.0131984010248522, -0.330624559129269, -0.178529511448759, 
    0.0410758729991616, -0.077797344743367, 0.134512154337116, 
    -0.218937700797494, -0.0137214460789446, -0.0604332454289641, 
    0.036048915625738, -0.252608499580276, -0.0199805352731218, 
    0.131132902630075, 0.141075362596928, 0.198068020502304, 
    0.24486837036872, 0.181518843684185, 0.160039367235615, 
    0.275519967688345, 0.307969463090243, 0.238001845730709, 
    0.19093345228693, 0.16775076360049, 0.157133463500686, 0.187726213335473, 
    0.22582354406831, 0.204438395277967, 0.186196117051962, 
    0.226113851314442, 0.229062759881729, 0.196667184599828, 
    0.203971906721898, 0.189277813686764, 0.15247062052203, 
    0.260268051968485, 0.28127142319182, 0.0997290631560509, 
    0.18935584111234, 0.527403020356669, 0.119667486165224, 
    -0.0527136937002883, -0.14289258507665, 0.624865083327473, 
    0.238155003187611, -0.124220380369957, 0.357111323772347, 
    0.466178219611786, 0.125433363576326, -0.208145818202214, 
    0.367094089063551, 0.542836416410594, 0.214910088263544, 
    -0.00995937601921708, -0.182628123093604, -0.171958279995629, 
    0.360709376734097, 0.217911273705939, 0.215443115444644, 
    -0.0175119844541015, 0.533962917229253, 0.0229804024750963, 
    -0.145517979757054, 0.0550828096782527, -0.117384791285847, 
    0.0399369976399943, -0.272449094411976, -0.00350852900496872, 
    -0.507416578944449, -0.208161279697457, -0.0529954940664184, 
    -0.310368712665717, -0.0674572145107524, 0.0888156612769935, 
    0.0894350876030017, 0.118042946339955, 0.0894543860751816, 
    0.0627544101706987, 0.148250950767929, 0.182816580605607, 
    0.122283088841239, -0.137332619103678, 0.238470932982538, 
    0.412705754563624, 0.162189967976763, 0.033937718105595, 
    -0.143284258383496, 0.190987267617778, 0.464798445665848, 
    0.381757957691873, 0.277302952311423, 0.194622451337833, 
    -0.104790440750941, 0.791574834854599, 0.275688425941473, 
    0.064417207656611, 0.239257141644447, -0.401109080334222, 
    0.492540963228999, 0.44292473418954, 0.201862536076418, 
    -0.139838682594963, 0.200356507870534, 0.384518887152963, 
    0.0273718329781497, -0.0706256109765629, -0.115635001972035, 
    0.00318104273482797, 0.446603663722809, 0.237190520667455, 
    0.037812127437776, 0.236765452906405, 0.149445155737084, 
    0.100441065214492, 0.414865151742592, 0.197331413632409, 
    -0.0056801247750382, 0.047618199102789, 0.314835182078304, 
    0.0971776550914158, -0.0234728495284664, 0.18181802300292, 
    0.191638273498356, 0.146673921651055, 0.018122715479228, 
    -0.0828751887088016, -0.0435874550337475, -0.0301381580943287, 
    -0.0105976311052652, -0.0752082532401438, 0.0109787292991105, 
    -0.0205851113353165, -0.148381057669289, -0.0157602897052402, 
    -0.127067313736498, 0.021931490510726, -0.155065837119625, 
    0.0101152093710335, -0.269385838667948, -0.10078443086078, 
    -0.023745455210842, -0.219181748429993, 0.0154757057841027, 
    0.0618708983696465, 0.0697443354200349, 0.108642881161398, 
    0.147749852409427, 0.134253927025601, 0.143129663663119, 
    0.194351547511844, 0.126973751498949, 0.0163798744412714, 
    0.350793288963452, 0.293192382328495, 0.0222721169021563, 
    0.047322538499227, 0.591021444888268, 0.336149975363202, 
    0.0964989035353548, 0.0183746921074856, 0.303199376460901, 
    0.322575876074417, 0.219038252674467, 0.608555498069861, 
    0.514895288284286, -0.00544368778213485, 0.555261316575399, 
    0.79767368247857, -0.137728450157445, -0.312675906284058, 
    0.274749345309048, 0.391879689292796, -0.108261799290083, 
    -0.0167758500006739, -0.0783435320548217, -0.0123171451082661, 
    0.0316861418723386, -0.0224938154158189, -0.0361199367216697, 
    -0.0430268501048559, 0.00581318033396516, -0.0122250345628266, 
    0.0717677197410835, 0.0817360940912354, 0.0783418694151648, 
    0.0810729371041405, 0.0738442546639275, 0.0736148028764733, 
    0.0737387595141315, 0.0769997018630985, 0.0270938747217524, 
    0.11235909933208, 0.273863853015222, 0.0708604138512099, 
    -0.0192937400037521, 0.344574245964541, 0.290989605178819, 
    0.129117495454191, 0.501652824079115, 0.355829973779225, 
    -0.160017512497894, 0.256648603929709, 0.513448416515201, 
    0.0724859073217662, 0.664618390572327, 0.64738595787211, 
    0.0134280276192086, 0.313915251356708, 0.852224458206944, 
    0.507256901298812, 0.262119652211181, 0.0816557751422823, 
    -0.125970471547747, 0.260958393452478, 0.319570746245694, 
    0.11070653581302, 0.280598198204455, 0.546022883954935, 0.22137005826233, 
    -0.0528767551601899, 0.234805834091511, 0.493335080685785, 
    0.159404194447983, 0.0694798721126572, -0.208087711680537, 
    0.445906264263266, 0.313871929029603, -0.0565519922288027, 
    0.425894979634114, 0.495242122209273, -0.0660451928663345, 
    -0.0321585177644471, -0.30194925472456, 0.25111355588629, 
    0.381627367134335, 0.171554494545341, 0.155171151140011, 
    0.529370900567475, 0.226410872553832, -0.221930134327042, 
    0.399608040384175, -0.12404172093739, -0.451128025015696, 
    -0.0228787319039033, -0.349894490413289, -0.038448694518439, 
    -0.297787894930286, 0.00622797886122083, -0.257412731708517, 
    0.0904261151640897, -0.303586956502998, 0.00697308473778407, 
    -0.0904904489502939, 0.111838334218541, 0.00739997295598076, 
    0.100973424970981, 0.024142092043304, 0.0975053924507174, 
    0.0164256774583443, 0.064717024204994, -0.182750880573171, 
    0.0159242676531803, -0.0463602585028751, -0.0337264821312279, 
    -0.0657320591565618, -0.0299199876126672, -0.0227232762297576, 
    -0.0537028487503939, -0.0116285816590151, 0.0126556620724795, 
    0.0108704983043092, -0.0604614308514602, 0.024382386860022, 
    0.00679931847653731, 0.00958105096349521, 0.0102828966143696, 
    0.00900557431419963, 0.00834924885641107, 0.0102567991190208, 
    0.0204010586586175, 0.0176171781140993, -0.146607475693641, 
    0.481503005487277, 0.106699666169943, -0.12214513082469, 
    -0.046049721480701, 0.34116838158197, 0.584053028899852, 
    0.301100430772694, 0.179431242662771, 0.605893049739456, 
    0.0981501006834582, -0.0144119227819759, -0.0721125701102805, 
    0.342615957740197, -0.0812251470501512, 0.166222721596242, 
    0.453838972058575, 1.22545078844436, 0.797704030388965, 
    -0.0278670742868017, -0.108717759669898, -0.168452340704095, 
    -0.0201992589388794, -0.125261770595038, -0.0800554801134643, 
    -0.100189707828631, -0.080247211936091, -0.0898061380290843, 
    -0.0665626648763184, -0.0606526227069527, -0.0495411625188139, 
    0.269515713104663, -0.0722235812338667, 0.21163316762715, 
    0.444463729552689, 0.211483251258886, 0.121700609207187, 
    -0.187818191381595, 0.334042411410425, 0.367372898103012, 
    0.153331455968037, -0.0676017049033333, 0.444597073425943, 
    0.265570147862401, 0.0161108546388186, -0.0246168387269397, 
    0.580530932769319, 0.20897666032831, -0.0670373235387187, 
    0.20797869384022, 0.435549609792358, 0.116403771824977, 
    0.059530672453803, 0.0655548918039987, 0.0644472188678614, 
    0.0673033041084198, 0.0703330691727955, 0.0771089461614683, 
    0.0640698393116473, 0.0407814982580878, 0.0406001756268383, 
    0.183038916633863, 0.062513917691009, 0.20395484162199, 
    0.333848280549718, 0.211187500905233, 0.205859934593584, 
    0.171273243972396, -0.0550993712251505, 0.398190614907096, 
    0.499553892239368,
  -0.0402300519737001, -0.541443062553906, 0.366522936864857, 
    0.396376296150815, -0.0845462091563854, -0.107408110173388, 
    0.267338350832905, 0.488405625980646, -0.0773759061611155, 
    0.864640214510529, 0.299851478764135, -0.0270080927751378, 
    -0.0460176878525763, -0.0584819464211529, -0.0327954443545494, 
    -0.17115192701308, -0.040050919526041, 0.0104351370415959, 
    -0.0723305525395555, 0.00228164059449235, 0.160828100395437, 
    0.123721031929893, 0.0778853371513915, -0.0147497346100082, 
    0.030759507250621, 0.200440551964063, 0.124539872420373, 
    0.0321959530260198, 0.0893111700166266, 0.135921399699875, 
    0.113101615296912, 0.121749050170601, 0.182570586105821, 
    0.171194210373177, 0.151687144614382, 0.164183875405616, 
    0.15474950573379, 0.154630253209094, 0.17910111567035, 0.188410469029418, 
    0.202201580721817, 0.192498654789488, 0.186344246286467, 
    0.206215214532937, 0.213446576085766, 0.176214153469781, 
    0.189587144855613, 0.266768590564931, 0.204691770523913, 
    0.167414535987935, 0.238764920448236, -0.167545328719977, 
    0.623510540899446, 0.439576998859988, 0.0133336793402895, 
    -0.0829296179654728, -0.248159460298403, 0.11835343197924, 
    0.788310778887818, 0.177249165923626, -0.0595628620750695, 
    0.0372148346575621, 0.0459666286959698, -0.0114581605975876, 
    0.887940398256467, 0.298765640547595, -0.132720508951925, 
    0.450964703848846, 0.386606653502134, -0.0145777864637831, 
    -0.169240895790204, 0.0735834146324687, -0.12748306175043, 
    0.0163321012224802, -0.244321544622325, -0.0464890478295394, 
    -0.120722365272856, -0.204329606580756, 0.211151141726743, 
    -0.126643748196223, 0.201634447014239, 0.0768331951897886, 
    0.168119462312296, 0.370827969881282, 0.117313364538858, 
    -0.158094850817586, 0.428667138027266, 0.724835287216798, 
    -0.0215591801324297, -0.547638440923762, -0.00763436341261828, 
    0.71299905427075, 0.00566512401737915, -0.00802862203723956, 
    0.205879704280986, -0.500125829040757, 0.645112352959187, 
    0.49893918760312, 0.049066237887183, 0.23191833180189, 0.577181827827169, 
    0.270684590435088, -0.0663937864738522, -0.0848206070969224, 
    -0.272505195113528, 0.223995622242098, 0.272331164863604, 
    -0.357606048588088, -0.230573765032884, -0.00968527180047973, 
    -0.165732276457476, -0.049357923248151, -0.197454527709877, 
    0.0507260201842099, -0.0241733070956099, -0.132976388998782, 
    0.0382196403392332, -0.123651893313782, -0.173095023838465, 
    -0.00144398613006299, -0.170203622596999, -0.0475026826768531, 
    -0.0640388008061171, -0.126404084028608, -0.0107364369804885, 
    -0.145954350756433, -0.10066165474736, -0.0221971535845697, 
    -0.045716165933723, -0.0186924447552233, 0.0945132031365607, 
    -0.153456970820308, 0.14992525116382, 0.322398278461912, 
    0.146402682054388, 0.0761540114282244, -0.146503862346942, 
    0.105569257773563, 0.207819234017045, 0.329443916912101, 
    0.409334549206032, 0.163813710797225, 0.164855173569272, 
    -0.384842766251106, 0.595269648219732, 0.460875657091994, 
    0.223953370542262, 0.138905642746385, 0.135151809050598, 
    -0.113177812044805, 0.413135608763831, 0.538861173215269, 
    0.177932120786289, 0.0840945392443616, 0.42775422424041, 
    0.375165034870025, 0.0926538957852514, -0.112136500057983, 
    0.00363642480860035, 0.267491304539819, 0.219228698371487, 
    0.127578326528854, -0.0485375262302264, 0.282398244157957, 
    0.156550344279082, 0.0410691244401006, 0.123914587224325, 
    0.221111269508344, -0.00890143900473286, 0.218781592395305, 
    0.336827299105145, 0.094299474827814, 0.0379412034675271, 
    -0.00141191814089155, 0.191915293574978, 0.132667359504267, 
    0.0317000950607757, 0.092908735663403, 0.237687043990966, 
    0.0483666916692601, -0.0249970137816737, -0.0332243540062695, 
    0.0383937560076782, -0.029587317238539, 0.0174944023752979, 
    -0.0803807432661072, -0.0131599393492204, -0.0200519991956367, 
    -0.033719126384967, 0.0339318787695822, -0.00970169147246386, 
    0.119502863380204, 0.2386628721629, 0.0717020793617007, 
    0.0767478196014765, 0.179639099046925, 0.328314596603712, 
    0.524934884110406, 0.0730821991317957, -0.518063506899077, 
    -0.119154830085514, 0.84265209817119, 0.119822618272324, 
    -0.246662103958884, 0.301384278614458, 0.75349553135711, 
    -0.146781270658914, 0.241234523199437, 0.974889886170641, 
    0.0278931291245892, -0.0834398283539285, -0.0720091073279332, 
    0.124680934352639, -0.0940279656223967, -0.019805124850283, 
    -0.135230342798718, 0.00590604745559418, 0.102475732517253, 
    -0.198786860630994, -0.131207006458343, -0.2695667831154, 
    0.0861291780482532, -0.212645448553737, 0.0435691498547179, 
    -0.11197123297123, 0.162516313081672, -0.138022680023937, 
    0.128220787227854, -0.259827121816025, -0.0237259232829129, 
    -0.070645008321645, 0.0370386878187276, -0.0516311275837356, 
    0.0438015570947904, -0.0130292945968625, 0.0346370633084024, 
    -0.0842059913400136, -0.01122843263567, -0.0678754914923691, 
    -0.0876259376038564, 0.0412176709535978, 0.0594552608411757, 
    0.0813726732624716, 0.10935432328342, 0.125728107667809, 
    0.122147776061565, 0.113654760873244, 0.125924738141636, 
    0.0989777038401107, 0.0421074227262756, 0.215416979829343, 
    0.229608166589237, 0.0960670404308085, 0.0857270849002737, 
    0.408795550610516, 0.282240485482505, 0.0416526612096388, 
    0.157597879115404, 0.52030336499544, 0.212553547142723, 
    -0.0481032088010171, 0.367299374083602, 0.414751574618444, 
    -0.0323436957129059, 0.380877102164554, 0.645826224046203, 
    -0.0195370807793818, -0.027770155217703, -0.206586609706038, 
    0.6286011368389, 0.21300581142215, 0.0388726488937634, 0.067619788313166, 
    -0.0627726157600499, 0.409356107738738, 0.302134685946827, 
    0.277932027484373, 0.691591560457358, 0.310713325686737, 
    0.0311905437921377, -0.0700220201714437, -0.175601631805797, 
    -0.0176333367041153, -0.0763306639649796, 0.11876118593598, 
    0.0657724197372815, 0.0281466788507638, 0.179744000781726, 
    -0.0296828875178671, -0.0895705354264134, -0.034058853880999, 
    -0.104191690245085, 0.0548874470801575, -0.0371501191251109, 
    0.0473103881308896, -0.262467349848724, 0.023463534567322, 
    -0.191167404001381, -0.0839381023620176, -0.108831653073637, 
    0.126291549727817, -0.0241582894955664, 0.306651443128017, 
    0.245612167472147, 0.0613326163159681, -0.0279675677798792, 
    0.0929250077093201, -0.201341138889535, 0.428015405813, 
    0.300126444365944, -0.162011452435738, 0.432706568750557, 
    0.748032993497109, 0.0934414754104854, -0.40292951514528, 
    0.0268958894598893, 0.956062097903133, 0.459004179254539, 
    0.0569807246705767, 0.516939811246534, 0.561620958867261, 
    0.500120245024296, 0.271667640485685, -0.226482724272226, 
    0.368159762628996, 0.311688512260352, -0.00827570216053018, 
    0.0238060707205516, 0.514756351350982, 0.273188331341612, 
    0.183106010025799, 0.365072565549015, 0.0202031282531508, 
    -0.0291354903734433, 0.0790096108695055, 0.113698604926493, 
    -0.0135098167347999, 0.381528626883004, 0.0445685096252038, 
    -0.0300443984124755, -0.0296861031167689, 0.0167511652175121, 
    -0.00991776676515131, -0.0159789475682347, 0.009849787508129, 
    0.00251051906223521, -0.0527635853081594, 0.0849605767839854, 
    0.0843697251868136, -0.102778553818177, -0.0186308340150781, 
    -0.0965476311954896, 0.418524625169759, 0.386273012019251, 
    0.168353765364737, 0.262067521260928, 0.337108313375443, 
    -0.229391328535005, 0.0292590375196571, 0.890312874051664,
  -0.0300904971008755, 0.00710098370641853, -0.0195480734309562, 
    -0.0303351002164331, 0.0699293097703422, -0.0152369248643155, 
    0.0420642405272784, 0.0114452283328858, 0.0510122535508429, 
    -0.0462579643621145, 0.0836091963756373, 0.0940439363505906, 
    0.0274032423762643, 0.274548315491885, 0.245626164935023, 
    0.0604484257918931, -0.0575994571063457, 0.0325568372568307, 
    0.458209919599087, 0.305379940712447, 0.0278104743404491, 
    0.515534183675522, 0.385600823767672, 0.0635093656360351, 
    -0.175676943602929, 0.049294755272312, 0.72256669884996, 
    0.172245514078001, -0.217205837997503, 0.258703216473415, 
    0.480242842264822, -0.155995489504953, -0.0962062395130165, 
    0.0428107859677042, -0.152696149415283, 0.00178115177320039, 
    0.177942233982811, -0.00630520616463193, -0.00705883859622641, 
    0.209526208225673, -0.0906032725852568, 0.122867282500171, 
    -0.202581460809799, 0.0538919015723752, -0.247437725266133, 
    -0.0157165110267594, -0.472572515305987, -0.150031222498125, 
    -0.119068009893469, -0.297742057478772, -0.153639364577121, 
    0.130741747107739, 0.137242003487231, 0.0360330762513657, 
    0.00471442079880551, 0.173020607683829, 0.320200905186194, 
    0.241483737988439, 0.080131509576827, 0.0539927903060467, 
    0.626668733164206, 0.263414779092744, -0.063749692661448, 
    -0.20151205646447, 0.746617856715623, 0.56797447711455, 
    0.178106933758523, 0.0795367858629249, -0.217275373437599, 
    0.931819042002392, 0.329595849384677, 0.0563823925351678, 
    -0.417611885120655, 0.249515452421081, 0.666461058683932, 
    0.169281431988819, 0.138225862368528, -0.267712212676712, 
    0.435252269121448, 0.226594174421856, -0.032557564446552, 
    0.0447391038076282, 0.367116719965126, -0.2463808220143, 
    0.0272797122427824, -0.286178462113433, 0.175652927248997, 
    -0.116550782933924, 0.220656468229611, -0.157707727030595, 
    -0.45077112855752, -0.06596683031683, -0.107616370907802, 
    0.174281020966835, -0.641663726720783, 0.0669445203186258, 
    -0.225460412003515, -0.121526829087327, 0.0197310924843932, 
    -0.583295495354321, -0.0856311460236877, 0.0332091519710853, 
    0.0888903437021466, 0.0560613267489316, 0.0279374573557903, 
    0.192610199447472, 0.244916892370037, 0.141994342201001, 
    0.0623488188085592, -0.0351924163392758, 0.302180560993358, 
    0.30626945114481, 0.160217307023818, 0.172505519159373, 
    0.259524571033627, 0.175471993797815, 0.414680291479631, 
    0.584194429491803, 0.293371995748997, 0.144183007464756, 
    -0.241389459692988, 0.529667268718727, 0.369106769901595, 
    -0.00760756176258622, 0.347936906761819, 0.627248960613678, 
    -0.0693609199788484, 0.0881243899624317, -0.330049724533968, 
    0.293773106171608, 0.462814667837678, 0.233693536505295, 
    -0.0159017250810796, 0.526339790457559, 0.410066870334382, 
    0.254817481466366, 0.278478406498079, 0.157870831674679, 
    -0.0954479009214461, -0.307012275474608, 0.221047074431499, 
    0.788061985922342, 0.0211411953091457, -0.207924532425216, 
    0.00682629798973648, 0.453621369536796, 0.0171301170110548, 
    0.221006255903732, 0.672510969766679, 0.153925413288667, 
    0.00322185387806775, -0.154814657687031, 0.0613013515440039, 
    0.356139898821969, 0.0726900658933331, -0.0198702040088654, 
    -0.0418489882727003, 0.223916843077231, 0.148982807115724, 
    0.0362060667565397, 0.202862477757048, 0.265163363153023, 
    0.099469985761852, -0.0116916185454578, 0.0533695486680862, 
    0.249631328649173, 0.150177168424054, 0.0455062761134481, 
    0.0529530923673624, 0.300611145554222, 0.263524861390317, 
    -0.135067864197156, 0.22862087866744, 0.47580084866823, 
    0.355336775165279, 0.173227277269849, -0.244008904820974, 
    0.0717902451793253, 0.358683037294678, 0.16978898871198, 
    0.311217140589325, 0.452024074099822, 0.0735727916443197, 
    -0.0224283235627165, 0.112199297540724, 0.352127181127715, 
    0.0144562166509606, 0.299887574387117, 0.442339657422004, 
    0.0279606550114751, -0.050769889715829, -0.0679558633725964, 
    0.0126885157972532, -0.0683698897953518, -0.0171583888677199, 
    -0.0716258944668421, -0.0363767543057927, -0.0254066934876254, 
    -0.0421563695062497, 0.00525855561912232, 0.13252916672571, 
    -0.0528786549050492, 0.267157516687114, 0.24342912317185, 
    0.0676729699446518, 0.0558626020595759, 0.219378897460745, 
    0.548705724792677, 0.0333694992980112, -0.343685840217604, 
    -0.182545590224727, 0.518890082224084, 0.14166273526547, 
    0.788105106527908, 0.944922343192784, 0.192918118112735, 
    -0.384956019947789, 0.465028092949471, 0.897690385392042, 
    -0.0810151898768418, -0.186328303423896, -0.084476888548133, 
    -0.119990681308986, -0.145264819462119, -0.0158832252423061, 
    -0.0868054461774594, -0.15378604816978, 0.0466080198989375, 
    -0.169692923026229, 0.0272944279276909, -0.121927491258112, 
    0.0181342259175093, -0.0739709554589002, 0.0354212634240247, 
    -0.108082836158537, 0.00953669097775019, -0.0913635503315901, 
    -0.0632598376703213, -0.00176898851690402, -0.0740940235805993, 
    -0.0270109334663004, 0.079040269275531, 0.171397285645517, 
    0.0962254392302204, 0.168515048605629, 0.338334111465495, 
    0.181204276470257, 0.023489631616027, 0.0627999640775409, 
    0.303384917378667, 0.289577522959104, 0.201489223887852, 
    0.158489586419292, 0.156191277795189, 0.16707016872044, 0.14805757909872, 
    0.105048360109965, 0.139522528362803, 0.241952913641148, 
    0.149417417368703, 0.0146549173916117, -0.000753385737059506, 
    0.0419024567546727, 0.0170994256554895, 0.0339269520470967, 
    0.0212405230177932, 0.0358333299460846, 0.0299619354111067, 
    0.0415254838802252, -0.0128758693390895, 0.0439880866173221, 
    0.0828385056079997, 0.119879292498815, 0.148383046005912, 
    0.141775786819116, 0.0990131987771883, 0.0677341429551808, 
    0.148256684635606, 0.204449308713763, 0.156322716416843, 
    0.347930750733893, 0.263129305164583, -0.303222261784748, 
    0.334925616289875, 0.429893622142903, 0.039513323828211, 
    0.474123339394982, 0.556212025645535, 0.17663144672717, 
    0.126229315436628, -0.196626116763209, 0.263584210718472, 
    0.127424294398527, 0.0790797875165394, 0.106718775606041, 
    -0.134937549849547, 0.182297605009414, 0.198014532631258, 
    0.0701372209006791, -0.0268378269183899, -0.102104577790651, 
    -0.139665898697645, 0.194031444914031, -0.343380841602913, 
    0.0927626271796657, -0.202809670188001, 0.100088581790156, 
    -0.174276651935945, 0.167272224229111, -0.221668569036836, 
    0.144020247685457, 0.0700100775593344, 0.0483328818780687, 
    0.0695738661661701, 0.095746518800125, 0.0933478729147042, 
    0.128524056476886, 0.155910526423752, 0.105236631071731, 
    0.048748768412253, 0.136762819040089, 0.158551514638962, 
    0.123918706565348, 0.214663688286639, 0.289936423536706, 
    0.143083960767772, 0.142036926389324, 0.45630609150538, 
    0.164819665410349, 0.0419203838229663, -0.142329099560592, 
    0.45957468385868, 0.319756860767836, 0.149382074197218, 
    0.104073726474853, 0.172451120139502, -0.171493291768708, 
    0.64717833493569, 0.41147436264866, 0.0574598764909078, 
    0.0522808688614672, 0.436849398137063, 0.307580546050799, 
    0.275675810962838, 0.182266427968968, -0.231056147118072, 
    0.103802413383947, 0.220705660920221, 0.45483680949189, 
    0.458470950388714, -0.0202578699466069, -0.111121437306493, 
    -0.109671104587076, -0.120882006905783, -0.16864355242409, 
    -0.134960991049486, -0.108148429111888, -0.149134997338523, 
    -0.0654608811932535, -0.162452637652055,
  0.159360232141321, 0.0134223963749163, 0.37843489539109, 0.518125351167363, 
    0.0308994385271204, -0.0944012863155372, -0.096816463796909, 
    0.544362911622664, 0.070356427376618, -0.203720052525487, 
    0.296175097085486, 0.273926077639009, 0.0989713868966318, 
    -0.252947348559911, 0.46943708088489, 0.286072131138009, 
    0.0922245026935369, 0.0990856569920658, 0.517518237947717, 
    0.0955914968938319, -0.0583749878921412, -0.0744047372451053, 
    0.0572862196078711, -0.0336295686703302, 0.0602693687878094, 
    -0.0746179054261057, 0.0396496692317835, -0.030955272708125, 
    0.0584077275363242, -0.105447579846178, 0.0273521272204667, 
    0.120267199409801, 0.157938271925433, 0.156591122506014, 
    0.178826487672861, 0.205354856551078, 0.240986299081063, 
    0.290125887021504, 0.225057342658173, 0.118485367958672, 
    0.258435262924714, 0.362534918515082, 0.293622427581157, 
    0.406120204966645, 0.371824967327426, 0.0494652967771154, 
    0.296611860026208, 0.613329769444907, 0.333309369607223, 
    0.508419843585826, 0.396851907541371, -0.255668118204245, 
    0.284701739153523, 0.528819265158313, 0.119780139634956, 
    -0.379435770437952, 0.657931946190314, 0.541003051115365, 
    0.226498362206572, 0.156072083887227, 0.140100388599581, 
    0.337537182913433, 0.163358583947427, -0.0492189876227749, 
    -0.131802036861446, -0.0217182587129045, 0.0899418773604065, 
    -0.0034965110391168, 0.197635144800482, 0.0921951734644503, 
    -0.0105196983037941, -3.83351650874858e-05, 0.000476685549036959, 
    0.00294439943040559, 0.00213480871403003, 0.0057368558270475, 
    -0.0228227838679696, 0.0664066605869915, 0.0835673544947282, 
    -0.147187370150625, 0.045267612281496, 0.263485045224302, 
    0.118789086692746, 0.306330217338062, 0.229636849021863, 
    0.0589428203975849, 0.637502967565013, 0.406969247667683, 
    0.000246592270872689, -0.244140335629557, 0.0403288400709928, 
    0.126070368996538, 0.175168791320173, 0.966866898346513, 
    0.836685563128652, 0.222013123254536, -0.671824729957569, 
    0.202179554838599, 0.651807406671114, 0.320449866243073, 
    0.168954389806748, 0.287997250499546, 0.13826911864372, 
    0.0591834562110908, 0.0411311772710018, 0.0346717615041593, 
    0.0385712950157885, 0.045022371334512, 0.0181413485755679, 
    0.0572657867480088, 0.186954928764071, 0.0312836001030559, 
    -0.0289589389009526, 0.340378886271615, 0.248921516469739, 
    0.120611315399824, -0.0498506951993274, 0.351497825754367, 
    0.179293817789816, -0.0906956340591727, 0.0694712211364522, 
    0.445499854765548, 0.387925593648476, 0.246807355352179, 
    0.152527816957974, 0.241222248595463, 0.21642457886814, 
    0.937067099425943, 0.222613810699384, -0.0582656899550711, 
    -0.124442117509581, -0.16025835532348, -0.0803103933165001, 
    -0.103417208023082, -0.125403458867595, -0.117757696021105, 
    -0.0758438238875218, -0.0956555666362386, -0.0654697575735829, 
    -0.120772014298683, 0.0537309769121895, 0.0135084066970545, 
    0.0647974098878227, 0.028811042805199, 0.0518889596023322, 
    -0.0320401125881485, 0.0296305014620549, -0.000239305890212912, 
    0.009246157726778, 0.0744845227844927, -0.00708294172092853, 
    0.15107490761824, 0.217814171423584, 0.182384567194444, 
    0.131751952218017, -0.102626918413793, 0.292774375874821, 
    0.237847426532515, -0.0459166234228187, -0.201936081692444, 
    0.27175129428327, 0.250114294745091, 0.0361345119579337, 
    -0.532402708835518, 0.28815227110339, 0.258778714502802, 
    0.656218302850162, 1.07129773844842, -0.171625583308083, 
    -0.307533979340958, -0.233958951786473, -0.0745099087687473, 
    -0.173679009857713, -0.127472439527538, -0.175433227308312, 
    -0.149582908426737, -0.12269893186522, -0.179816334138955, 
    -0.0409528574861804, -0.166331497888362, 0.0525479865774066, 
    0.0614042357873249, 0.113797382244666, 0.0424048732340967, 
    0.0712877232109595, 0.137284293780001, 0.156540599589064, 
    0.122182666665497, 0.126751978705079, 0.0156571606904456, 
    -0.00773625319568974, -0.116331172293472, 0.00945968919209736, 
    -0.0743914116259272, -0.0138061121338759, -0.0234918858462685, 
    0.0358776485590272, -0.0583883110605915, 0.0547986979392496, 
    -0.135132264930655, -0.000827886449072779, 0.0123481119559266, 
    0.0531209852106963, 0.0574737106418647, 0.0442764354260348, 
    0.0394052799532542, -0.0879692307453312, 0.288215134678435, 
    0.0968229807542252, -0.327911037029138, 0.0365418861633932, 
    0.466505880950916, 0.0789307760432226, -0.24289741059893, 
    0.495126024768361, 0.541056145558328, 0.0747283036252866, 
    -0.0530463544814786, -0.0899482447267236, 0.241361500536361, 
    0.133639499529849, 0.281610814009283, 0.527860382695863, 
    0.355327193139985, 0.106360810053533, 0.244635461881409, 
    0.657799885014207, -0.0555614867584495, -0.242586197095867, 
    0.0518015938715594, -0.309296935890544, -0.152657497966545, 
    -0.130764452520379, -0.233729560656264, 0.0144475087814535, 
    -0.215991090539906, 0.0594168262620312, -0.170487818280746, 
    0.0693959327292469, -0.234838871411161, -0.0125200588981192, 
    0.077301073336693, 0.0816034101202056, 0.125079233550058, 
    0.176881580014059, 0.17484306313395, 0.207544291847233, 
    0.158432813208988, -0.0861949023619991, 0.363270592561124, 
    0.39408923599484, 0.0190309277127441, -0.0530542546572738, 
    0.600521070825426, 0.371042909041369, 0.14552489930238, 
    -0.0299210283143821, -0.0704932173580246, -0.0356924449355538, 
    0.770883073143588, 0.272676746696645, -0.242022687815801, 
    -0.195017923159655, -0.488052173376646, 0.143302157292791, 
    0.651261127504815, -0.00625451038732985, -0.37133504016044, 
    0.0477015607819082, 0.427999188237882, 0.000388394111527121, 
    0.00852817108064202, -0.116102217366609, 0.00369344221327196, 
    -0.18813450665072, -0.0349175032402101, -0.217143305374817, 
    -0.138049686215901, -0.00444478392363901, -0.191423488499244, 
    0.0275520994707114, 0.0228680045744104, 0.263229312897407, 
    0.328956635677336, 0.143491590228941, -0.178707464587166, 
    0.345365442307817, 0.466732665041371, 0.0628126551886559, 
    -0.0544776797841863, 0.167197526187589, -0.193705542024108, 
    0.137007059861873, 0.996408040773576, 0.154305778994992, 
    -0.159648878959845, 0.122094110722429, 0.282701473708576, 
    0.340290726706212, 0.711657823621859, 0.46775620276172, 
    0.413599839676191, 0.530855972331154, 0.228086847215909, 
    0.0470540083698039, -0.369578721063085, 0.234155729012846, 
    -0.0309560655630417, -0.0873142428041857, -0.0901523424750362, 
    -0.0608678161413868, -0.444176579097355, 0.173974692831777, 
    -0.126191049014093, 0.0698347992779908, -0.0994539593931424, 
    0.0894182712603998, -0.181978498674935, 0.0741349141238907, 
    -0.112434518698104, 0.178104380598141, -0.0995179228758988, 
    -0.0136236022662011, 0.00980037204398855, 0.0602562236924959, 
    0.0230513557620895, 0.0973510738379515, 0.064274257819458, 
    0.0674902475501351, 0.0346858784166787, 0.233581769778432, 
    0.12623056487648, 0.0237072261073396, 0.165697778742145, 
    0.283749158853014, 0.230037726409572, 0.167962846794243, 
    0.0955331367586161, 0.0690850601174722, -0.296410501694281, 
    0.515981524224942, 0.373137158472415, -0.125797306010371, 
    0.36462472246543, 0.581573684082533, 0.291654249545408, 
    0.151768514631157, -0.308691660382702, 0.151212006229658, 
    0.540552004647109, 0.223407237731691, 0.110063863523788, 
    0.0703029890837686, 0.12801601332007, 0.160657719793046, 
    0.183932305165088, 0.409835956737835, 0.440501333673364, 
    0.237950381636441, 0.139779789656753,
  0.939667727473292, -0.211916522998552, -0.0516825324204712, 
    -0.211190800808912, 0.269575452802785, 0.554734773726777, 
    0.132736119318213, -0.305439552182147, 0.269258550922825, 
    0.538027276995845, -0.419755000604563, -0.116062438203004, 
    -0.227840817395804, -0.0895924386709612, -0.23085118845765, 
    -0.083683693195561, -0.200547449469263, -0.208596485950063, 
    -0.0475030673874738, -0.231738599018202, 0.0375781006263914, 
    0.00548501216243663, 0.19083815327012, 0.192846338137407, 
    0.116554276655213, 0.0978522982701641, 0.135505995486812, 
    0.124530816443782, 0.0415619697907255, 0.0621185904088575, 
    0.122551999607051, 0.12629285521484, 0.0998432037198776, 
    0.0786187764694911, 0.0689492319901664, 0.0802671900944479, 
    0.074349546407025, 0.0660136003670942, 0.0574331600287612, 
    0.0755594805190176, 0.0535648933541072, 0.0754541687956942, 
    0.0621870291073887, 0.0497377858403204, 0.080121052685942, 
    0.0712933189866799, 0.0815134478294198, 0.0895073707946506, 
    0.0835381929175578, 0.0503760542033619, 0.120751744177532, 
    0.0804976965975958, 0.125734669837439, 0.291357563741325, 
    0.196457611162217, 0.030944032330379, 0.105240563081286, 
    0.44079514586902, 0.0954496847801484, -0.0876459900476501, 
    -0.133731035775838, 0.140761786338576, 0.585866488127574, 
    0.468427905912459, 0.0585932407592096, -0.102031510204195, 
    -0.280901056312565, 0.282767345906726, 0.522904804129947, 
    0.210351537022962, 0.0158721687540671, 0.149899836067989, 
    -0.111980901869413, 0.233281363615778, 0.2560165286671, 
    0.115560479672684, 0.368430426028058, 0.237407335727999, 
    -0.00627649120255706, -0.0573693146312403, -0.0900050794201997, 
    -0.195764339168089, 0.0510362502995906, -0.0830988688337603, 
    0.0517918113956328, -0.159455380649997, 0.0454911691249966, 
    -0.155213907196333, 0.00511874619668033, -0.184063523776967, 
    -0.0448040827727309, 0.0370486807246324, 0.203625662123175, 
    0.167597843175061, 0.0423287049602048, 0.0113689197865523, 
    0.399818710365693, 0.27140321217651, 0.155056344040666, 
    -0.422971393661818, 0.282790336903918, 0.563988713089007, 
    0.157182796484803, 0.0562078828500459, -0.264049273882339, 
    0.561468382703693, 0.325946289036848, 0.145834831919983, 
    -0.125417814131665, 0.371231045007684, 0.303776809548791, 
    0.20508523014544, 0.0974216060955893, -0.0369406166701321, 
    -0.121689833094655, 0.194384294339895, 0.379205336076357, 
    0.0626542706775055, -0.0218339358630611, 0.0946809884988834, 
    -0.215177545013322, 0.0983745894821175, -0.355476713754671, 
    -0.043692754206815, -0.221514052916326, -0.21373797249813, 
    0.0517343745648292, -0.167242211578852, 0.138678479597074, 
    -0.155363835075712, 0.12266241013273, -0.0154443213345045, 
    0.0270479484382975, 0.0211598253160763, 0.0532775260768335, 
    0.0134200057399387, 0.0578893413365606, 0.00753588191127799, 
    0.0315249716613574, -0.0600748429623746, -0.000479105216803305, 
    0.0645053056921286, 0.0703814178532195, 0.0574228214457067, 
    0.0751278654147541, 0.0726823658784115, 0.139035287943393, 
    0.163935429346284, -0.0169424420241752, 0.0388654493028708, 
    -0.338504541445324, 0.171960553819724, 0.492554890391539, 
    0.207034556120284, -0.0700721870417111, 0.0151782901186831, 
    0.32667521208411, 0.655007670838986, 0.310405351788719, 
    0.025233431686493, 0.0174172982554346, 0.370334557934757, 
    0.0892020224604928, 0.0419127105536297, -0.0127194965390845, 
    0.206442035764582, 0.468054363622575, -0.130505710767443, 
    -0.105304929742944, -0.111772263857604, -0.456433178947381, 
    -0.196614769830658, 0.0224445105037044, -0.161315974103846, 
    0.267835094010097, -0.436190815419915, 0.0772843875849502, 
    -0.367689100860228, -0.134575993776594, -0.177067526074206, 
    -0.0451823515073607, 0.110836545909991, 0.0599681713105368, 
    0.048866096649247, 0.0439999089341691, 0.10020870584163, 
    0.156786184981572, 0.0920622597805509, 0.0115478984052323, 
    0.0521618871045519, 0.0813976530082557, 0.0917825860287463, 
    0.0966428979495927, 0.119373496947572, 0.134140598068999, 
    0.0873007703818244, 0.079089485274298, 0.29040418556324, 
    0.017606302288722, -0.0742051574558633, -0.101164341304547, 
    0.470889039437119, 0.16254543950838, -0.0266080481855211, 
    -0.244560971231504, 0.467826799526208, 0.697032831854596, 
    0.369501759704514, 0.031946715066011, -0.312548597759099, 
    -0.150675405007251, 0.240210290596074, 0.215285418929239, 
    0.786090751158534, 0.516497974570195, 0.0361889806550788, 
    0.0938646891976157, 0.798643490723092, 0.020336762928018, 
    -0.0582493643481155, -0.266806076271218, -0.175188824929092, 
    0.0276369337651398, -0.13811485821552, 0.0831822302236293, 
    -0.238724111011193, -0.0648968715467417, -0.0631364611349457, 
    -0.0796759510946784, -0.0995670660060514, -0.243916928221942, 
    0.197828495821145, 0.294171072473417, 0.0792632265941727, 
    0.00406220572715524, -0.0938191498761114, 0.515049297505456, 
    0.116660022138044, 0.0979882262993449, -0.191240267086595, 
    0.569302690478185, 0.327609512225987, 0.0724054685987144, 
    -0.203922043535722, -0.283994687016255, 0.456311285557039, 
    0.674556645712471, 0.204344294605029, -0.221521739918046, 
    0.153717169547664, 0.514963685570185, 0.138750664944503, 
    -0.159263205440444, 0.237518218154044, 0.375117406889889, 
    0.0241591903623291, -0.151692765323086, -0.0348782484521963, 
    0.413483353653065, 0.143802246020987, 0.0508519046260622, 
    0.0746142030272854, -0.122391964425706, 0.435863415253001, 
    0.198825409628157, 0.0617446944384615, -0.137381788374764, 
    0.061006092053545, 0.233217969765953, 0.251542541141349, 
    0.282967501685329, 0.23055200080604, 0.105840006857799, 
    0.0341414036995062, -0.0200035750307416, -0.0872609861850695, 
    -0.0305646151888791, 0.351535670103394, 0.15919175547555, 
    0.0171130828580384, -0.0379499382928129, 0.102891441256071, 
    -0.139847796433847, 0.00115437673362687, -0.340318514161617, 
    -0.137287917491422, -0.0253930625728673, -0.184065741460561, 
    -6.43738125593041e-05, -0.182481853496423, -0.0350667494927368, 
    0.0619353864183594, 0.120619263048991, 0.0692779147254753, 
    0.0815303971015956, 0.274251778281857, 0.255840232411944, 
    0.0769380627462067, 0.0800583808288717, -0.359546272868751, 
    0.506633149558303, 0.361810542694041, 0.242558820876323, 
    0.763452521029102, 0.240069455740672, 0.105991778473016, 
    -0.391547737164524, 0.473278154982183, 0.552884311562758, 
    0.127587388907345, -0.152098306317716, -0.0569233056142819, 
    0.31164883002242, 0.236812009743884, 0.315991567112159, 
    0.484571373690842, 0.0424160163947608, -0.312216559217044, 
    0.00149532461632221, 0.417858428068087, -0.0795650565454766, 
    -0.16183470028461, -0.254149477220906, -0.286547565235476, 
    -0.127094464291382, -0.158703019777681, -0.133956993895446, 
    -0.042896798854575, -0.142523890706955, -0.0493719016363765, 
    -0.059035852022298, 0.248427031454256, -0.175288999262576, 
    0.0696373907241443, -0.0238259590023789, 0.0814409590905299, 
    -0.356830523032421, 0.0115442571724946, -0.326576874984472, 
    -0.280754105247224, -0.0142081317061913, -0.0323306724185151, 
    -0.04680872733249, 0.0539354773394271, -0.0267028980723162, 
    -0.067382834099976, -0.0457851656905382, -0.0863007525772474, 
    0.183992789131884, 0.0546642409329565, -0.228933640124473, 
    0.104489028431012, 0.64643514993136, 0.0530029025100523, 
    0.0427081943090968, 0.965208035734646, 0.268960863632291, 
    0.0760963003801455, 0.108044653372331, -0.0848229420054249,
  -0.0408906636604045, -0.110730591956218, 1.12506409970972, 
    0.00051514467143722, -0.442101136925877, 0.0201951017882824, 
    0.969734287735437, 0.228856362991154, 0.0308980996952601, 
    0.00487796734824784, 0.330042793685197, 0.257876134666813, 
    0.162121726299246, 0.0973796303261664, -0.0298332696145958, 
    -0.288397150622171, 0.0731279751793897, 0.293939654352663, 
    -0.244209209247349, -0.177703683355745, -0.0355584080082617, 
    -0.297764965820992, -0.0550461198819506, -0.170557621071708, 
    -0.213911654477143, 0.0417025468540508, -0.171791551683935, 
    0.0894308033576227, -0.219820805517211, 0.00457519443051006, 
    -0.00646086763312472, 0.0819612817106091, -0.012670088563797, 
    0.0786185923377145, -0.0322047182116008, 0.0717787879332805, 
    -0.0343159699195215, 0.0562191465249294, -0.0721034760751381, 
    0.00680451351329837, -0.0453313639557825, -0.0638378309135936, 
    0.0303943207783207, -0.00571283864932989, 0.0441360791739958, 
    -0.0375653615049755, 0.04164135528443, -0.015207027403294, 
    0.130851044363568, -0.106720032589579, 0.171855733913684, 
    0.214700614026685, 0.123376149004328, 0.0839677631079402, 
    -0.114368751467034, 0.22620368693101, 0.468136157474625, 
    0.0493288574713884, 0.00507613543297958, -0.134483407535942, 
    0.558881536010141, 0.19360741782446, 0.0746767747376625, 
    -0.118305173749915, -0.116141899600206, 0.0196473213672795, 
    0.644860188357552, 0.654183231365825, 0.12818539995317, 
    -0.149382067864257, -0.0494538593018135, 0.46013009716805, 
    0.291184296118499, 0.213765045317625, 0.240486222899486, 
    0.14225815003439, -0.24740155222555, 0.49708266666177, 0.325339705913833, 
    -0.000122765516004528, 0.751333675609063, 0.47801677379416, 
    -0.0116673891380581, -0.0845781306719078, -0.188946050513316, 
    0.549873572203858, 0.263447871249779, 0.11321794726478, 
    -0.164751998439517, 0.142932065179657, 0.100101794526178, 
    0.222172647034647, 0.756318415875237, 0.348557441152374, 
    0.137364878728388, -0.038777177340558, 0.700342895598121, 
    -0.0701246265615356, -0.312406918672762, 0.160638093779568, 
    0.354479761830612, -0.0250982191229787, -0.0604104385600568, 
    0.0573641782215078, 0.0724872712885597, -0.0196509942043642, 
    0.0760728232544284, 0.0912863917103073, -0.000301146614367975, 
    -0.0729661984977988, 0.148111324820135, 0.162042690889243, 
    -0.0318497957058399, 0.0463015334518639, 0.306650484743938, 
    0.168340933707787, 0.0454493766765736, 0.26836623931794, 
    0.265637455061166, -0.0540286198522382, 0.482723815026414, 
    0.313173886878794, -0.00119804714323546, 0.212544721453113, 
    0.464780404352293, 0.0511281429559606, -0.115088234730159, 
    0.218861256609935, 0.258126968472395, 0.0171945083188899, 
    -0.0728347676807913, -0.173185666459623, 0.0793195009011193, 
    -0.153805324592353, 0.0189349968812843, -0.28373598814044, 
    -0.101898796697927, -0.042056630069388, -0.201890680254636, 
    0.0415867608548447, -0.0358413371341788, 0.0592128512015055, 
    0.00651582697277334, 0.0369816107918336, 0.0397245948925665, 
    0.0452095273462658, -0.0302737589260716, 0.0263260356688306, 
    -0.0558897226557513, -0.04702946780005, 0.0412916924745399, 
    0.0361438826958113, 0.0398153394430448, 0.0378559484583858, 
    0.0342530427313049, 0.034410679620626, 0.0371010159269796, 
    0.0547212339961663, 0.0732673373855224, -0.014051642287117, 
    0.0134273381591776, 0.183857859659959, 0.245033198765511, 
    0.15514473016691, 0.0926012108160937, 0.0401104160429468, 
    0.181460772650024, 0.595349391098121, 0.0892875665630504, 
    -0.340435461564818, 0.140822860637701, 0.556161855674228, 
    -0.0051299220735431, -0.136834299180161, 0.346929720169195, 
    0.764196304504521, -0.346036992800023, -0.451001329699463, 
    0.612383720119407, -0.427634943632943, -0.49963730641434, 
    -0.161336549141826, -0.074258629534759, -0.219109801995387, 
    0.0113443810295666, -0.263539168946407, -0.0435354896902001, 
    -0.419796063809263, -0.0701502114772898, -0.389935549962176, 
    -0.0420537009252557, -0.257655327227043, -0.0975256393085892, 
    -0.116852716967741, -0.0676878828748659, -0.430816895631596, 
    0.0104233058561748, -0.0770838332580194, 0.0523760848958374, 
    -0.283604664350565, -0.0731578550414056, 0.118341885692952, 
    0.0914697386155017, 0.0286898010021723, 0.125249368706967, 
    0.198119328537917, 0.113267171064078, 0.0629228525783064, 
    0.130387320741073, 0.183257218993739, 0.199188176152859, 
    0.164022467969995, 0.192315948628833, 0.210846772087808, 
    0.181245821840811, 0.172823905978149, 0.162314180110159, 
    0.163755919128864, 0.142206603168702, 0.161260970732937, 
    0.33058483794125, 0.218851191396678, 0.0452343661679707, 
    0.0162947422604456, 0.367723151733118, 0.34116589951234, 
    0.130345624010082, -0.0688025089191164, 0.066571470298755, 
    0.41759003982563, 0.29700389399931, 0.0438865732738684, 
    -0.0372290715036862, 0.150640567445777, 0.86864018620783, 
    0.389961674113307, -0.0583028727781619, 0.235184756502568, 
    0.7114053685588, 0.224718215921204, -0.203326543819057, 
    0.136227573380699, 0.791240170425755, 0.339044048534428, 
    -0.211797038089387, 0.577281482543129, 0.38050797089165, 
    -0.0612618453161941, 0.322827565655758, 0.613281920174559, 
    0.159290368139818, 0.057948471516305, -0.0407841928881885, 
    0.12405934352605, -0.190638130987455, 0.165285373070061, 
    0.338754470542227, -0.0237021525652394, -0.0668876920703298, 
    -0.0193454377499816, 0.213896732183706, 0.1041358484753, 
    0.0843123758523206, -0.0400235207967224, 0.0903642971803763, 
    0.184901624234576, 0.138212968441607, 0.0749542696379868, 
    -0.101986287128424, 0.275294350234699, 0.236767453760319, 
    0.00147176254857093, -0.143226271450768, 0.226998765448877, 
    0.460641162552144, 0.211530776765791, -0.137123981548838, 
    0.271861388844272, 0.397485589540166, 0.104324621531414, 
    -0.0138091891332028, -0.0728635724708525, 0.440530782100577, 
    0.203838676156718, 0.0171272535283034, 0.102520893465286, 
    0.367803169642904, 0.129539383571976, -0.0829400515632112, 
    0.151658714750811, 0.371710165447425, 0.261357258128829, 
    0.156578623917371, 0.144691907076005, 0.190392710968994, 
    0.130678457369486, 0.0479743129091615, 0.269911370939184, 
    0.129480545400242, -0.0267994837790776, -0.103211945436729, 
    0.41946629947376, 0.324974067671584, 0.221527115616718, 
    -0.202750383512725, 0.540148519669403, 0.29308686193615, 
    -0.0881926430973669, 0.293360558634309, 0.413137170053375, 
    0.250223205566212, 0.929126030465604, 0.404131484032746, 
    0.0877749220135691, 0.16500550591086, -0.00234159189226589, 
    0.686335242992912, 0.213707810039607, 0.220012624023445, 
    0.173742499611073, -0.317673711140367, -0.323112588583007, 
    -0.125970869216553, -0.275495607133179, -0.123030914364431, 
    -0.292367226517983, -0.152970075618558, -0.0554613304195577, 
    -0.273996357900759, -0.0248659980725012, -0.0336815374422188, 
    0.155840629003182, 0.0078822081181253, 0.0206287653313709, 
    -0.158483977070728, -0.0551252529967983, 0.0547503765088533, 
    0.0172123671413976, 0.131853424149859, -0.0264770541126855, 
    0.0378731076886011, -0.0694033283992948, -0.0249458157020621, 
    -0.0232446460405157, -0.0103322591302063, -0.0355063970189622, 
    -0.0387867933419735, 0.0236162272366927, -0.00838481393055919, 
    -0.0370025102302274, -0.103670340825925, 0.0277786539222319, 
    0.282108094627856, 0.156528924644984, 0.0337869249033486, 
    0.200724926319524, 0.290399088547913, -0.111119640619355, 
    0.360562130230573, 0.320266906040724,
  0.547497927059475, 0.141327496452566, -0.0216528554846673, 
    -0.0709670153043605, 0.0302798602710198, 0.115735361024181, 
    -0.104795530489107, 0.0523913546446246, 0.205057151284903, 
    -0.0253916679891889, 0.0354667619432031, 0.0222097939852895, 
    0.392956997165495, 0.0971617857989696, 0.0185852123142966, 
    0.139206261097976, 0.242705119707403, -0.0242950878793667, 
    0.0208769170380065, 0.385713050249861, 0.38228086055024, 0.2267638101612, 
    -0.0671870104482383, 0.498714384688014, 0.201105815036581, 
    0.0727381555768482, -0.333956961341423, 0.396681110671444, 
    0.435426280523039, 0.109413931581434, -0.0963866376990646, 
    0.0437708738110655, -0.13585148542633, -0.0258385741167695, 
    -0.100645801273959, -0.0580984512407373, -0.0715512574642088, 
    -0.0743607185930139, -0.0135507443827381, -0.0978991448845774, 
    0.0300821812470743, 0.0717172877616705, 0.128616594393212, 
    0.152422813940601, 0.122620257395119, 0.153659371786334, 
    0.244808704846285, 0.157678256917615, -0.0171168148612157, 
    0.207988419901539, 0.429577588128782, -0.0350183510893936, 
    0.105613502693223, 0.649105457133024, 0.40823935470752, 
    0.085889605026276, -0.0696169070318081, -0.226475447744319, 
    0.624282606275772, 0.122917249514826, -0.118859810114354, 
    0.186374698523627, 0.450500172613319, 0.00157396483613871, 
    0.48991973061956, 0.43093616110323, 0.222756207293259, 0.919124444302329, 
    0.518646616696575, 0.0268186091804253, -0.0925128180074387, 
    0.0471176730904852, -0.176465703109901, -0.0445010098067959, 
    -0.073155284656949, -0.108909583071425, -0.0116741085551675, 
    -0.0243315920472618, 0.0696055183926582, -0.143689502052563, 
    0.112543625986746, 0.138545649914818, -0.0173471784171727, 
    0.317821221928813, 0.484365660680931, 0.156784308380661, 
    -0.247482998947575, 0.237140421272027, 0.612444990025892, 
    0.137975155872046, -0.397857110799281, 0.347769021456298, 
    0.519548869999074, -0.00983348757853381, 0.184961679353778, 
    -0.386801924092289, 0.540968800694408, 0.480565417586714, 
    0.204600976192663, -0.187844942155341, 0.029682880932133, 
    0.442872283071131, 0.311464718973988, 0.166432749693421, 
    0.072293102107791, 0.0649498759657065, -0.333702331149055, 
    0.359046853870342, 0.337618288775862, 0.22705258743809, 
    0.343152030050913, 0.143365435293479, -0.0348059638993001, 
    0.286396380720687, 0.030290735533028, -0.129740824886839, 
    0.00636415352011731, 0.290133670911662, -0.118398205732371, 
    -0.0472294286390834, -0.0182319175106972, -0.224895206890632, 
    0.102105697224982, -0.0386503462453624, 0.0752504672013574, 
    -0.158256932804005, 0.0365980957658405, -0.0847946561126418, 
    0.0387425751286869, -0.227667206063906, -0.0367589424107387, 
    0.114351751806881, 0.155823349065099, 0.136018943772345, 
    0.164758252576915, 0.197479711707039, 0.190217568386756, 
    0.210904354023469, 0.321706143692408, 0.444433726410555, 
    0.301861537558016, 0.0383856271127973, -0.0995337105586346, 
    0.760780764896812, 0.434408217189727, 0.110276808594521, 
    -0.154476320994251, 0.747157104086888, 0.374310717591575, 
    0.0855577203669829, -0.178988047429227, 0.556185930552677, 
    0.389755603182545, 0.0534171016670824, -0.0865606540481585, 
    -0.171586595725672, 0.430134996656645, 0.462870693625486, 
    0.139458796601445, -0.246991032085546, 0.171360770253786, 
    0.387102352883223, 0.144954076192315, 0.122509855059227, 
    -0.239894618713511, 0.271576728548234, 0.31241192400801, 
    0.0957083699537394, -0.018203738317445, 0.0576244894501894, 
    0.143046132177413, 0.338471759002515, 0.195019474267921, 
    0.0384882555327068, 0.0603459363483852, -0.137521772699252, 
    0.0938010273045117, 0.104704032610311, 0.245435287576286, 
    0.159019036749568, -0.0165675989647122, 0.0328478691205041, 
    -0.231239688885307, -0.0081070979813502, -0.205485463690791, 
    -0.195678227390072, 0.0457288394532791, -0.0589025291094521, 
    0.10551476125525, -0.171682112229358, 0.0373330411089586, 
    0.0767878267845493, 0.0768104841617249, 0.107108952724387, 
    0.114901997466371, 0.0863299018689854, 0.0927220781688597, 
    0.128796480817926, 0.10919964238725, 0.0563750488476326, 
    0.107207043055355, 0.127609082065438, 0.167116340700263, 
    0.252627105707278, 0.321409772258786, 0.203833412818907, 
    0.00213343909803446, 0.113610151591094, 0.531352009391404, 
    0.191698732935166, 0.0211471077113611, 0.253425887067, 0.399241218139103, 
    0.00583447321230711, -0.258130511358703, 0.286261216889773, 
    0.706511892925311, 0.386069480181108, 0.324344715676153, 
    0.616791245383854, 0.245665844131135, 0.0579489907903356, 
    0.0163320364537727, 0.0170422900507367, -0.0964188232487927, 
    0.0492398713218498, 0.0953196229081267, -0.277152895411523, 
    -0.166335028755909, -0.138071253866863, -0.0834965740118508, 
    -0.226598787805303, 0.104579754091845, -0.113097590067173, 
    0.117517005405323, -0.159552519826681, 0.0292388303890231, 
    -0.0571972895258869, 0.066505540518101, -0.251127528281364, 
    0.0164033976650814, 0.050622811382266, 0.0708399067092638, 
    0.073487884998018, 0.0758314707458615, 0.0422340984090562, 
    0.0518073594490984, 0.0868609009169215, 0.0646357923763774, 
    0.00105087628542465, 0.0726868905506342, 0.102594820208252, 
    0.214621778109716, 0.195280617371926, 0.0210666010039579, 
    0.242143364769865, 0.351719304422933, 0.011239595565957, 
    -0.0200826893023687, -0.0771437202386909, 0.410900280363622, 
    0.112346033836721, 0.630652780180086, 0.48163200136672, 
    -0.0428328574461888, 0.0900502463213922, 0.168090328672822, 
    -0.398642326376328, 0.138579171792012, 0.604089257390911, 
    0.122398512751494, 0.0936619736299482, 0.217165017067217, 
    0.00206258664472175, -0.0745883340677015, -0.0920213387562182, 
    0.0105235111586817, -0.15365521992566, 0.0035688500205618, 
    0.00501976806943752, -0.172305224168264, 0.109140960594203, 
    -0.299239423375336, -0.0309149493054587, -0.164969883833818, 
    -0.223674158111434, 0.0964177350502161, -0.135955107969684, 
    0.0572100630169093, -0.239953407561425, -0.0177324364961606, 
    0.0206619917697395, 0.070405365926775, 0.134518439939407, 
    0.119789329635996, 0.0663181341687991, -0.126319081803735, 
    0.43341173810314, 0.305010235792828, -0.104318238013255, 
    0.611091186261233, 0.301194964806663, 0.00942484832072296, 
    -0.0763681808190872, 0.737489612035313, 0.393182945119882, 
    0.147242588227868, -0.227330506654647, -0.129373463124219, 
    0.667884808136494, 0.130361308797713, -0.0375292026796074, 
    -0.214283087540436, -0.0627822358029441, 0.821134056034386, 
    0.339223735407879, 0.287438237585724, 0.320816685022948, 
    -0.333986106282076, 0.00045507400410412, -0.340187676985156, 
    0.0217434438695913, -0.305049242966522, -0.190740568248303, 
    -0.106447806321934, -0.229019117962462, -0.0206433621488802, 
    -0.209064564282227, 0.0286320805560107, -0.23747494736924, 
    -0.0264036074091351, 0.117839469300046, 0.101453085388341, 
    0.0875699397156332, 0.161098524407272, 0.240545913320404, 
    0.329708235899395, 0.168143419877331, -0.166994397354809, 
    0.149926015862794, 0.475387189913705, 0.101147857529982, 
    0.538476519845136, 0.647130670142423, 0.219314174906643, 
    0.14095736815341, -0.118169503730987, 0.722233226436124, 
    0.47557710316067, 0.212556283266326, -0.0667470062459609, 
    -0.0527197061595466, -0.00134750865817662, 0.986180439323333, 
    0.325178821081407, 0.00600557800499667, -0.104983703256484, 
    0.131889943683488, 0.185815430665689, 0.640857425276997 ;


 X_priorinf_mean = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 X_priorinf_sd = 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 Y_priorinf_mean = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
                   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 Y_priorinf_sd = 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6,
                 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 time = 1000.0 ;

 advance_to_time = 1000.0 ;

}

