netcdf perfect_input {
dimensions:
	member = 1 ;
	metadatalength = 32 ;
	location = 960 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;

	double state(time, member, location) ;
		state:long_name = "the model state" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

// global attributes:
		:title = "true state from control" ;
                :version = "$Id$" ;
		:model = "Lorenz_04" ;
		:model_scale = "2-scale" ;
		:model_forcing = 15. ;
		:model_delta_t = 0.001 ;
		:space_time_scale = 10. ;
		:coupling = 3. ;
		:K = 32 ;
		:smooth_steps = 12 ;
		:time_step_days = 0 ;
		:time_step_seconds = 3600 ;
		:history = "same values as in perfect_ics r813 (circa July 2004)" ;
data:

 MemberMetadata =
  "true state" ;

 location = 0, 0.00104166666666667, 0.00208333333333333, 0.003125,
    0.00416666666666667, 0.00520833333333333, 0.00625, 0.00729166666666667,
    0.00833333333333333, 0.009375, 0.0104166666666667, 0.0114583333333333,
    0.0125, 0.0135416666666667, 0.0145833333333333, 0.015625,
    0.0166666666666667, 0.0177083333333333, 0.01875, 0.0197916666666667,
    0.0208333333333333, 0.021875, 0.0229166666666667, 0.0239583333333333,
    0.025, 0.0260416666666667, 0.0270833333333333, 0.028125,
    0.0291666666666667, 0.0302083333333333, 0.03125, 0.0322916666666667,
    0.0333333333333333, 0.034375, 0.0354166666666667, 0.0364583333333333,
    0.0375, 0.0385416666666667, 0.0395833333333333, 0.040625,
    0.0416666666666667, 0.0427083333333333, 0.04375, 0.0447916666666667,
    0.0458333333333333, 0.046875, 0.0479166666666667, 0.0489583333333333,
    0.05, 0.0510416666666667, 0.0520833333333333, 0.053125,
    0.0541666666666667, 0.0552083333333333, 0.05625, 0.0572916666666667,
    0.0583333333333333, 0.059375, 0.0604166666666667, 0.0614583333333333,
    0.0625, 0.0635416666666667, 0.0645833333333333, 0.065625,
    0.0666666666666667, 0.0677083333333333, 0.06875, 0.0697916666666667,
    0.0708333333333333, 0.071875, 0.0729166666666667, 0.0739583333333333,
    0.075, 0.0760416666666667, 0.0770833333333333, 0.078125,
    0.0791666666666667, 0.0802083333333333, 0.08125, 0.0822916666666667,
    0.0833333333333333, 0.084375, 0.0854166666666667, 0.0864583333333333,
    0.0875, 0.0885416666666667, 0.0895833333333333, 0.090625,
    0.0916666666666667, 0.0927083333333333, 0.09375, 0.0947916666666667,
    0.0958333333333333, 0.096875, 0.0979166666666667, 0.0989583333333333,
    0.1, 0.101041666666667, 0.102083333333333, 0.103125, 0.104166666666667,
    0.105208333333333, 0.10625, 0.107291666666667, 0.108333333333333,
    0.109375, 0.110416666666667, 0.111458333333333, 0.1125,
    0.113541666666667, 0.114583333333333, 0.115625, 0.116666666666667,
    0.117708333333333, 0.11875, 0.119791666666667, 0.120833333333333,
    0.121875, 0.122916666666667, 0.123958333333333, 0.125, 0.126041666666667,
    0.127083333333333, 0.128125, 0.129166666666667, 0.130208333333333,
    0.13125, 0.132291666666667, 0.133333333333333, 0.134375,
    0.135416666666667, 0.136458333333333, 0.1375, 0.138541666666667,
    0.139583333333333, 0.140625, 0.141666666666667, 0.142708333333333,
    0.14375, 0.144791666666667, 0.145833333333333, 0.146875,
    0.147916666666667, 0.148958333333333, 0.15, 0.151041666666667,
    0.152083333333333, 0.153125, 0.154166666666667, 0.155208333333333,
    0.15625, 0.157291666666667, 0.158333333333333, 0.159375,
    0.160416666666667, 0.161458333333333, 0.1625, 0.163541666666667,
    0.164583333333333, 0.165625, 0.166666666666667, 0.167708333333333,
    0.16875, 0.169791666666667, 0.170833333333333, 0.171875,
    0.172916666666667, 0.173958333333333, 0.175, 0.176041666666667,
    0.177083333333333, 0.178125, 0.179166666666667, 0.180208333333333,
    0.18125, 0.182291666666667, 0.183333333333333, 0.184375,
    0.185416666666667, 0.186458333333333, 0.1875, 0.188541666666667,
    0.189583333333333, 0.190625, 0.191666666666667, 0.192708333333333,
    0.19375, 0.194791666666667, 0.195833333333333, 0.196875,
    0.197916666666667, 0.198958333333333, 0.2, 0.201041666666667,
    0.202083333333333, 0.203125, 0.204166666666667, 0.205208333333333,
    0.20625, 0.207291666666667, 0.208333333333333, 0.209375,
    0.210416666666667, 0.211458333333333, 0.2125, 0.213541666666667,
    0.214583333333333, 0.215625, 0.216666666666667, 0.217708333333333,
    0.21875, 0.219791666666667, 0.220833333333333, 0.221875,
    0.222916666666667, 0.223958333333333, 0.225, 0.226041666666667,
    0.227083333333333, 0.228125, 0.229166666666667, 0.230208333333333,
    0.23125, 0.232291666666667, 0.233333333333333, 0.234375,
    0.235416666666667, 0.236458333333333, 0.2375, 0.238541666666667,
    0.239583333333333, 0.240625, 0.241666666666667, 0.242708333333333,
    0.24375, 0.244791666666667, 0.245833333333333, 0.246875,
    0.247916666666667, 0.248958333333333, 0.25, 0.251041666666667,
    0.252083333333333, 0.253125, 0.254166666666667, 0.255208333333333,
    0.25625, 0.257291666666667, 0.258333333333333, 0.259375,
    0.260416666666667, 0.261458333333333, 0.2625, 0.263541666666667,
    0.264583333333333, 0.265625, 0.266666666666667, 0.267708333333333,
    0.26875, 0.269791666666667, 0.270833333333333, 0.271875,
    0.272916666666667, 0.273958333333333, 0.275, 0.276041666666667,
    0.277083333333333, 0.278125, 0.279166666666667, 0.280208333333333,
    0.28125, 0.282291666666667, 0.283333333333333, 0.284375,
    0.285416666666667, 0.286458333333333, 0.2875, 0.288541666666667,
    0.289583333333333, 0.290625, 0.291666666666667, 0.292708333333333,
    0.29375, 0.294791666666667, 0.295833333333333, 0.296875,
    0.297916666666667, 0.298958333333333, 0.3, 0.301041666666667,
    0.302083333333333, 0.303125, 0.304166666666667, 0.305208333333333,
    0.30625, 0.307291666666667, 0.308333333333333, 0.309375,
    0.310416666666667, 0.311458333333333, 0.3125, 0.313541666666667,
    0.314583333333333, 0.315625, 0.316666666666667, 0.317708333333333,
    0.31875, 0.319791666666667, 0.320833333333333, 0.321875,
    0.322916666666667, 0.323958333333333, 0.325, 0.326041666666667,
    0.327083333333333, 0.328125, 0.329166666666667, 0.330208333333333,
    0.33125, 0.332291666666667, 0.333333333333333, 0.334375,
    0.335416666666667, 0.336458333333333, 0.3375, 0.338541666666667,
    0.339583333333333, 0.340625, 0.341666666666667, 0.342708333333333,
    0.34375, 0.344791666666667, 0.345833333333333, 0.346875,
    0.347916666666667, 0.348958333333333, 0.35, 0.351041666666667,
    0.352083333333333, 0.353125, 0.354166666666667, 0.355208333333333,
    0.35625, 0.357291666666667, 0.358333333333333, 0.359375,
    0.360416666666667, 0.361458333333333, 0.3625, 0.363541666666667,
    0.364583333333333, 0.365625, 0.366666666666667, 0.367708333333333,
    0.36875, 0.369791666666667, 0.370833333333333, 0.371875,
    0.372916666666667, 0.373958333333333, 0.375, 0.376041666666667,
    0.377083333333333, 0.378125, 0.379166666666667, 0.380208333333333,
    0.38125, 0.382291666666667, 0.383333333333333, 0.384375,
    0.385416666666667, 0.386458333333333, 0.3875, 0.388541666666667,
    0.389583333333333, 0.390625, 0.391666666666667, 0.392708333333333,
    0.39375, 0.394791666666667, 0.395833333333333, 0.396875,
    0.397916666666667, 0.398958333333333, 0.4, 0.401041666666667,
    0.402083333333333, 0.403125, 0.404166666666667, 0.405208333333333,
    0.40625, 0.407291666666667, 0.408333333333333, 0.409375,
    0.410416666666667, 0.411458333333333, 0.4125, 0.413541666666667,
    0.414583333333333, 0.415625, 0.416666666666667, 0.417708333333333,
    0.41875, 0.419791666666667, 0.420833333333333, 0.421875,
    0.422916666666667, 0.423958333333333, 0.425, 0.426041666666667,
    0.427083333333333, 0.428125, 0.429166666666667, 0.430208333333333,
    0.43125, 0.432291666666667, 0.433333333333333, 0.434375,
    0.435416666666667, 0.436458333333333, 0.4375, 0.438541666666667,
    0.439583333333333, 0.440625, 0.441666666666667, 0.442708333333333,
    0.44375, 0.444791666666667, 0.445833333333333, 0.446875,
    0.447916666666667, 0.448958333333333, 0.45, 0.451041666666667,
    0.452083333333333, 0.453125, 0.454166666666667, 0.455208333333333,
    0.45625, 0.457291666666667, 0.458333333333333, 0.459375,
    0.460416666666667, 0.461458333333333, 0.4625, 0.463541666666667,
    0.464583333333333, 0.465625, 0.466666666666667, 0.467708333333333,
    0.46875, 0.469791666666667, 0.470833333333333, 0.471875,
    0.472916666666667, 0.473958333333333, 0.475, 0.476041666666667,
    0.477083333333333, 0.478125, 0.479166666666667, 0.480208333333333,
    0.48125, 0.482291666666667, 0.483333333333333, 0.484375,
    0.485416666666667, 0.486458333333333, 0.4875, 0.488541666666667,
    0.489583333333333, 0.490625, 0.491666666666667, 0.492708333333333,
    0.49375, 0.494791666666667, 0.495833333333333, 0.496875,
    0.497916666666667, 0.498958333333333, 0.5, 0.501041666666667,
    0.502083333333333, 0.503125, 0.504166666666667, 0.505208333333333,
    0.50625, 0.507291666666667, 0.508333333333333, 0.509375,
    0.510416666666667, 0.511458333333333, 0.5125, 0.513541666666667,
    0.514583333333333, 0.515625, 0.516666666666667, 0.517708333333333,
    0.51875, 0.519791666666667, 0.520833333333333, 0.521875,
    0.522916666666667, 0.523958333333333, 0.525, 0.526041666666667,
    0.527083333333333, 0.528125, 0.529166666666667, 0.530208333333333,
    0.53125, 0.532291666666667, 0.533333333333333, 0.534375,
    0.535416666666667, 0.536458333333333, 0.5375, 0.538541666666667,
    0.539583333333333, 0.540625, 0.541666666666667, 0.542708333333333,
    0.54375, 0.544791666666667, 0.545833333333333, 0.546875,
    0.547916666666667, 0.548958333333333, 0.55, 0.551041666666667,
    0.552083333333333, 0.553125, 0.554166666666667, 0.555208333333333,
    0.55625, 0.557291666666667, 0.558333333333333, 0.559375,
    0.560416666666667, 0.561458333333333, 0.5625, 0.563541666666667,
    0.564583333333333, 0.565625, 0.566666666666667, 0.567708333333333,
    0.56875, 0.569791666666667, 0.570833333333333, 0.571875,
    0.572916666666667, 0.573958333333333, 0.575, 0.576041666666667,
    0.577083333333333, 0.578125, 0.579166666666667, 0.580208333333333,
    0.58125, 0.582291666666667, 0.583333333333333, 0.584375,
    0.585416666666667, 0.586458333333333, 0.5875, 0.588541666666667,
    0.589583333333333, 0.590625, 0.591666666666667, 0.592708333333333,
    0.59375, 0.594791666666667, 0.595833333333333, 0.596875,
    0.597916666666667, 0.598958333333333, 0.6, 0.601041666666667,
    0.602083333333333, 0.603125, 0.604166666666667, 0.605208333333333,
    0.60625, 0.607291666666667, 0.608333333333333, 0.609375,
    0.610416666666667, 0.611458333333333, 0.6125, 0.613541666666667,
    0.614583333333333, 0.615625, 0.616666666666667, 0.617708333333333,
    0.61875, 0.619791666666667, 0.620833333333333, 0.621875,
    0.622916666666667, 0.623958333333333, 0.625, 0.626041666666667,
    0.627083333333333, 0.628125, 0.629166666666667, 0.630208333333333,
    0.63125, 0.632291666666667, 0.633333333333333, 0.634375,
    0.635416666666667, 0.636458333333333, 0.6375, 0.638541666666667,
    0.639583333333333, 0.640625, 0.641666666666667, 0.642708333333333,
    0.64375, 0.644791666666667, 0.645833333333333, 0.646875,
    0.647916666666667, 0.648958333333333, 0.65, 0.651041666666667,
    0.652083333333333, 0.653125, 0.654166666666667, 0.655208333333333,
    0.65625, 0.657291666666667, 0.658333333333333, 0.659375,
    0.660416666666667, 0.661458333333333, 0.6625, 0.663541666666667,
    0.664583333333333, 0.665625, 0.666666666666667, 0.667708333333333,
    0.66875, 0.669791666666667, 0.670833333333333, 0.671875,
    0.672916666666667, 0.673958333333333, 0.675, 0.676041666666667,
    0.677083333333333, 0.678125, 0.679166666666667, 0.680208333333333,
    0.68125, 0.682291666666667, 0.683333333333333, 0.684375,
    0.685416666666667, 0.686458333333333, 0.6875, 0.688541666666667,
    0.689583333333333, 0.690625, 0.691666666666667, 0.692708333333333,
    0.69375, 0.694791666666667, 0.695833333333333, 0.696875,
    0.697916666666667, 0.698958333333333, 0.7, 0.701041666666667,
    0.702083333333333, 0.703125, 0.704166666666667, 0.705208333333333,
    0.70625, 0.707291666666667, 0.708333333333333, 0.709375,
    0.710416666666667, 0.711458333333333, 0.7125, 0.713541666666667,
    0.714583333333333, 0.715625, 0.716666666666667, 0.717708333333333,
    0.71875, 0.719791666666667, 0.720833333333333, 0.721875,
    0.722916666666667, 0.723958333333333, 0.725, 0.726041666666667,
    0.727083333333333, 0.728125, 0.729166666666667, 0.730208333333333,
    0.73125, 0.732291666666667, 0.733333333333333, 0.734375,
    0.735416666666667, 0.736458333333333, 0.7375, 0.738541666666667,
    0.739583333333333, 0.740625, 0.741666666666667, 0.742708333333333,
    0.74375, 0.744791666666667, 0.745833333333333, 0.746875,
    0.747916666666667, 0.748958333333333, 0.75, 0.751041666666667,
    0.752083333333333, 0.753125, 0.754166666666667, 0.755208333333333,
    0.75625, 0.757291666666667, 0.758333333333333, 0.759375,
    0.760416666666667, 0.761458333333333, 0.7625, 0.763541666666667,
    0.764583333333333, 0.765625, 0.766666666666667, 0.767708333333333,
    0.76875, 0.769791666666667, 0.770833333333333, 0.771875,
    0.772916666666667, 0.773958333333333, 0.775, 0.776041666666667,
    0.777083333333333, 0.778125, 0.779166666666667, 0.780208333333333,
    0.78125, 0.782291666666667, 0.783333333333333, 0.784375,
    0.785416666666667, 0.786458333333333, 0.7875, 0.788541666666667,
    0.789583333333333, 0.790625, 0.791666666666667, 0.792708333333333,
    0.79375, 0.794791666666667, 0.795833333333333, 0.796875,
    0.797916666666667, 0.798958333333333, 0.8, 0.801041666666667,
    0.802083333333333, 0.803125, 0.804166666666667, 0.805208333333333,
    0.80625, 0.807291666666667, 0.808333333333333, 0.809375,
    0.810416666666667, 0.811458333333333, 0.8125, 0.813541666666667,
    0.814583333333333, 0.815625, 0.816666666666667, 0.817708333333333,
    0.81875, 0.819791666666667, 0.820833333333333, 0.821875,
    0.822916666666667, 0.823958333333333, 0.825, 0.826041666666667,
    0.827083333333333, 0.828125, 0.829166666666667, 0.830208333333333,
    0.83125, 0.832291666666667, 0.833333333333333, 0.834375,
    0.835416666666667, 0.836458333333333, 0.8375, 0.838541666666667,
    0.839583333333333, 0.840625, 0.841666666666667, 0.842708333333333,
    0.84375, 0.844791666666667, 0.845833333333333, 0.846875,
    0.847916666666667, 0.848958333333333, 0.85, 0.851041666666667,
    0.852083333333333, 0.853125, 0.854166666666667, 0.855208333333333,
    0.85625, 0.857291666666667, 0.858333333333333, 0.859375,
    0.860416666666667, 0.861458333333333, 0.8625, 0.863541666666667,
    0.864583333333333, 0.865625, 0.866666666666667, 0.867708333333333,
    0.86875, 0.869791666666667, 0.870833333333333, 0.871875,
    0.872916666666667, 0.873958333333333, 0.875, 0.876041666666667,
    0.877083333333333, 0.878125, 0.879166666666667, 0.880208333333333,
    0.88125, 0.882291666666667, 0.883333333333333, 0.884375,
    0.885416666666667, 0.886458333333333, 0.8875, 0.888541666666667,
    0.889583333333333, 0.890625, 0.891666666666667, 0.892708333333333,
    0.89375, 0.894791666666667, 0.895833333333333, 0.896875,
    0.897916666666667, 0.898958333333333, 0.9, 0.901041666666667,
    0.902083333333333, 0.903125, 0.904166666666667, 0.905208333333333,
    0.90625, 0.907291666666667, 0.908333333333333, 0.909375,
    0.910416666666667, 0.911458333333333, 0.9125, 0.913541666666667,
    0.914583333333333, 0.915625, 0.916666666666667, 0.917708333333333,
    0.91875, 0.919791666666667, 0.920833333333333, 0.921875,
    0.922916666666667, 0.923958333333333, 0.925, 0.926041666666667,
    0.927083333333333, 0.928125, 0.929166666666667, 0.930208333333333,
    0.93125, 0.932291666666667, 0.933333333333333, 0.934375,
    0.935416666666667, 0.936458333333333, 0.9375, 0.938541666666667,
    0.939583333333333, 0.940625, 0.941666666666667, 0.942708333333333,
    0.94375, 0.944791666666667, 0.945833333333333, 0.946875,
    0.947916666666667, 0.948958333333333, 0.95, 0.951041666666667,
    0.952083333333333, 0.953125, 0.954166666666667, 0.955208333333333,
    0.95625, 0.957291666666667, 0.958333333333333, 0.959375,
    0.960416666666667, 0.961458333333333, 0.9625, 0.963541666666667,
    0.964583333333333, 0.965625, 0.966666666666667, 0.967708333333333,
    0.96875, 0.969791666666667, 0.970833333333333, 0.971875,
    0.972916666666667, 0.973958333333333, 0.975, 0.976041666666667,
    0.977083333333333, 0.978125, 0.979166666666667, 0.980208333333333,
    0.98125, 0.982291666666667, 0.983333333333333, 0.984375,
    0.985416666666667, 0.986458333333333, 0.9875, 0.988541666666667,
    0.989583333333333, 0.990625, 0.991666666666667, 0.992708333333333,
    0.99375, 0.994791666666667, 0.995833333333333, 0.996875,
    0.997916666666667, 0.998958333333333 ;

 state =
   2.80267244662739,       2.56399157698841,       2.32223040073350,
   2.09702631702843,       1.86803760619422,       1.68039126579594,
   1.45791873297819,       1.32417405204412,       1.11597404368497,
   1.03234978914176,      0.857565484413053,      0.802573104400711,
  0.663866847629354,      0.633960253207987,      0.527951503475694,
  0.525319150791900,      0.449510972515386,      0.470177522695715,
  0.423845806889691,      0.459082597982086,      0.447290433081766,
  0.489580523784434,      0.513830906823197,      0.563644356369813,
  0.612592736544435,      0.671439114869410,      0.732687284221475,
  0.798346941454478,      0.865326518152282,      0.934191136309312,
   1.00286070339390,       1.07142077783311,       1.13865425672269,
   1.20444623752093,       1.26839733516248,       1.33054456815989,
   1.39108298002674,       1.45044160852948,       1.50918207860238,
   1.56816407472955,       1.62834203888589,       1.69125344782172,
   1.75786704752691,       1.83015780269364,       1.90902860005318,
   1.99648789286129,       2.09322274931047,       2.20100108645332,
   2.31973505389718,       2.45157147324842,       2.59831217796395,
   2.75955567169785,       2.93412931189614,       3.12162468922610,
   3.32147282999598,       3.53361059159070,       3.75621517937657,
   3.98905169318198,       4.23064601668987,       4.47951499252503,
   4.76052891494382,       5.02146816950991,       5.26525352692150,
   5.53625298593222,       5.82379289795485,       6.11993311984654,
   6.43173725893325,       6.74713352332771,       7.06664437699032,
   7.41070963753521,       7.77347065810400,       8.13545259323974,
   8.50257478743943,       8.88553191123127,       9.28468920379092,
   9.69718062661456,       10.1183667245061,       10.5448398172357,
   10.9763735371515,       11.4120743814158,       11.8462658592235,
   12.2734117178778,       12.6877637502539,       13.0796133598794,
   13.4580794241642,       13.8310440613846,       14.1531764212323,
   14.3996693736977,       14.6139267662445,       14.8143823822311,
   14.9670501887058,       15.0360860900786,       15.0155611734778,
   14.9161578526070,       14.8254321015701,       14.6794783659190,
   14.2014437925841,       13.7036386889489,       13.4070844570009,
   13.1955982568181,       12.6677960857503,       12.0582781041418,
   11.4825616469425,       10.9036083582878,       10.2907302486597,
   9.74612118010679,       9.22648704580800,       8.73437686621198,
   8.28723044040127,       7.73480988462400,       7.30465517271256,
   6.99972999702434,       6.54787606425494,       6.10320272736109,
   5.66135776393283,       5.19392173319898,       4.86483619671813,
   4.56382570655707,       4.10380357004102,       3.67528342757253,
   3.34205476892783,       2.91356293608774,       2.47077168761626,
   1.96873332112827,       1.60446525199815,       1.07426109657707,
  0.686343813821696,      0.151067258224355,     -0.247918193564739,
 -0.777996686059483,      -1.29241045909160,      -1.88721144522900,
  -2.22898375983363,      -2.89851843090804,      -2.80258239870343,
  -3.59292017662445,      -3.05218320509014,      -4.32010308782047,
  -2.92133865376036,      -3.74608237527841,      -3.13699218723905,
  -4.17186274866975,      -3.29448210780093,      -3.25418991217294,
  -2.58806091373469,      -3.47267547485786,      -2.45993608197491,
  -3.57438305108655,      -1.23359588450300,      -2.01954479389288,
  -1.40903057829824,     -0.782846657667618,     -0.204239984372007,
   1.10259636888402,       1.73688582456284,       2.74101866068023,
   3.47494935842845,       4.61532708352437,       5.24657577245537,
   5.95933817682820,       7.55387694360877,       8.40454740824460,
   8.55433618141343,       9.53829025538963,       10.3811217429337,
   9.66098000092698,       10.6790938650811,       10.9847784892026,
   9.67760260048162,       9.70646904692029,       10.8595362218513,
   10.6139277794878,       9.23277298515031,       8.96613045725664,
   8.50160000338879,       8.49964252842581,       7.33245075626003,
   6.78225640863553,       6.14600758002460,       5.32520490789616,
   4.71420116341202,       4.00267010313878,       3.61738850801983,
   2.95631283073549,       2.77513624250102,       2.21346198476345,
   2.16917475340367,       1.86689811184014,       1.89107881141505,
   1.83900305601990,       1.91962335037827,       2.05799060721310,
   2.24551485373150,       2.42517146854759,       2.61415753343859,
   2.73997837728296,       2.79805183385172,       2.86728304626652,
   2.89307906697999,       2.81524421548780,       2.71120218708209,
   2.57257664529016,       2.34223499004365,       2.05377927003863,
   1.74088930258490,       1.37198285072385,      0.973917121555087,
  0.555148403759069,      0.136112470227254,     -0.273568685996083,
 -0.679362688835729,      -1.05341526431974,      -1.30361366827495,
  -1.89485822019194,      -1.44629282636556,      -2.23411905486672,
  -1.67616499179950,      -1.96996092683687,      -1.88984903199036,
  -2.26584867865818,      -1.48373901910070,      -2.00566290971461,
  -1.49476014634351,      -1.65056198235066,      -1.37627053464542,
  -1.03683466019224,     -0.701284541837342,     -0.357676296727698,
  -2.36175742816489E-002, 0.439974344871406,      0.763551041144097,
   1.18185323093772,       1.55768870571512,       1.84063312773069,
   2.18016307362453,       2.49520495567557,       2.83406427597909,
   3.12166279698085,       3.24146979379452,       3.40984126516997,
   3.63290044099637,       3.84438796375237,       3.68569498259174,
   3.66888429927742,       3.70177648692110,       3.73556239568122,
   3.70990711211799,       3.52561678727919,       3.31179060355710,
   3.16087875750915,       3.03123295335190,       2.85341796755637,
   2.72055506331945,       2.54723508844817,       2.39366130553569,
   2.24835162721861,       2.19202753307682,       2.08484854223531,
   2.12435186277922,       2.10320214742005,       2.21603803581668,
   2.33169987390601,       2.50612848212889,       2.78688768465023,
   3.04944593406536,       3.46242318515870,       3.85243756324540,
   4.35147836857639,       4.87090845200504,       5.44792501281852,
   6.06161071755884,       6.70789276235145,       7.37958902405735,
   8.06743179897024,       8.76107865322486,       9.45209336250745,
   10.1309059482698,       10.7902430167137,       11.4180295425656,
   12.0029409053823,       12.5371499728255,       13.0184624762301,
   13.4440271436366,       13.8020025868240,       14.0809011849943,
   14.2873468336539,       14.4359892403137,       14.5245647854728,
   14.5329422298268,       14.4561853414894,       14.3145641924215,
   14.1234844298076,       13.8828357042293,       13.5767383728557,
   13.1856623762111,       12.7196218208718,       12.2059284792505,
   11.6533824275081,       11.0536034556210,       10.3990576244500,
   9.69590892988408,       8.95795319257722,       8.19428381888007,
   7.40978967303575,       6.60960219257803,       5.79957115253806,
   4.98640196784322,       4.17756517045648,       3.37988937590770,
   2.59897158321522,       1.83944206966745,       1.10522377285980,
  0.399463066175360,     -0.275721592716034,     -0.919354732100925,
  -1.53146194958875,      -2.11306269346381,      -2.66607814678129,
  -3.19324653510517,      -3.69801343231135,      -4.18435752341311,
  -4.65677560886161,      -5.12019323154001,      -5.57933266371374,
  -6.03782025091421,      -6.49759428925383,      -6.95853860173802,
  -7.41919206747297,      -7.87781321323636,      -8.33228136841750,
  -8.77976682295811,      -9.21687288084120,      -9.63971899904493,
  -10.0440042058738,      -10.4252215590950,      -10.7787441776766,
  -11.0999331939983,      -11.3842465021225,      -11.6273333493155,
  -11.8251302967274,      -11.9738762115680,      -12.0701648484928,
  -12.1110133317962,      -12.0939811144538,      -12.0172244870947,
  -11.8795564403866,      -11.6804290484860,      -11.4201211538029,
  -11.0996136213533,      -10.7206882065796,      -10.2859593725480,
  -9.79871116419873,      -9.26306669750643,      -8.68378961028868,
  -8.06634317876772,      -7.41667748517657,      -6.74128034490344,
  -6.04696431933620,      -5.34088160422741,      -4.63022850625406,
  -3.92232699390203,      -3.22432376079535,      -2.54317978297685,
  -1.88548135444585,      -1.25736886485558,     -0.664479497333985,
 -0.111836102995499,      0.396101212482811,      0.855475432049662,
   1.26307237352881,       1.61636770471762,       1.91351809229256,
   2.15339699496105,       2.33564871224960,       2.46070562697723,
   2.52978585688086,       2.54488557697491,       2.50877009833317,
   2.42493720726371,       2.29755074968469,       2.13136524050496,
   1.93163281239306,       1.70398985368703,       1.45434643589513,
   1.18876798436555,      0.913349393976909,      0.634103485039176,
  0.356840473304271,       8.70497496892113E-002, -0.170203822241739,
 -0.410380164513703,     -0.629533952758249,     -0.824377005291219,
 -0.992340602075095,      -1.13162946881414,      -1.24122471123994,
  -1.32085802913754,      -1.37098779965550,      -1.39275287158768,
  -1.38793222932975,      -1.35886625398606,      -1.30842539754107,
  -1.23994273934910,      -1.15699839116359,      -1.06314111840348,
 -0.961631900786283,     -0.855349560444707,     -0.747084732815463,
 -0.639116791781164,     -0.533379783240326,     -0.430728256026385,
 -0.331886863468612,     -0.236804651164188,     -0.145188998199419,
  -5.58650394278634E-002,  3.19319827764492E-002, 0.121233827359324,
  0.210722752769170,      0.308469793727750,      0.406925053193123,
  0.521731856940931,      0.638201453139567,      0.776439840961847,
  0.919982939294858,       1.08609615977724,       1.26332636864582,
   1.46083860261624,       1.67316644572430,       1.90279777255982,
   2.14774020779115,       2.40728622365126,       2.67889244011753,
   2.95982901880457,       3.24788592036895,       3.54235752993863,
   3.84056690287469,       4.13563875636676,       4.42172155710183,
   4.70065639169352,       4.97421035661078,       5.23453667419158,
   5.47279534919701,       5.68999500057107,       5.89705679097373,
   6.10345994937175,       6.28427649247657,       6.41516050117166,
   6.52157900406989,       6.63841537232636,       6.77743542205035,
   6.86003235410806,       6.88023231222867,       6.90553323652687,
   6.95265827090339,       7.03169086419997,       7.05478380277191,
   7.02268457778128,       7.02321605668267,       7.05295171078600,
   7.06497360770867,       7.05797456545607,       7.06400694439212,
   7.08018116300024,       7.10461137951073,       7.11792135193478,
   7.16380075935396,       7.19683589279064,       7.26587323458699,
   7.31920157406662,       7.39396524642080,       7.47389123553805,
   7.56236580368220,       7.65433772174020,       7.74787767658667,
   7.84529286813169,       7.94202745228966,       8.03336177335945,
   8.11666388510794,       8.18721144371567,       8.24403531477746,
   8.28531778810338,       8.30904282972873,       8.31136752077426,
   8.29195667515364,       8.25624214573935,       8.19590458968780,
   8.09097475876244,       7.95050153003047,       7.79693087542083,
   7.62940797776753,       7.43473916295147,       7.21222739531714,
   6.97062794827178,       6.71477844167965,       6.44291284503907,
   6.15849177740414,       5.86548258072551,       5.56301244198918,
   5.25440960467452,       4.94268156777633,       4.62686207290755,
   4.31074178123377,       3.99830948276134,       3.68746909532184,
   3.37876537661613,       3.07651324438306,       2.78101860721375,
   2.49200782198021,       2.21160743660234,       1.93984624502512,
   1.67576818588587,       1.42163754935909,       1.17961891854215,
  0.947475401737094,      0.723262792878788,      0.510605145142274,
  0.312195768413168,      0.123107443227391,      -6.08588400138922E-002,
 -0.234936308937261,     -0.394371455286016,     -0.544152528358034,
 -0.696201198815454,     -0.850486200987517,     -0.994747962896020,
  -1.12046418237910,      -1.24932574264713,      -1.40947615730366,
  -1.55853830405991,      -1.68029593901547,      -1.81183818617448,
  -2.00280273977221,      -2.15559515014000,      -2.30149963914586,
  -2.41960516560311,      -2.61057038319777,      -2.78837382577678,
  -2.92842688315299,      -3.07911115811900,      -3.24056031102335,
  -3.41124138405446,      -3.55438576943902,      -3.70945363887068,
  -3.85398727718000,      -3.99226815220500,      -4.12439491409212,
  -4.24747635992815,      -4.36116045541627,      -4.46772120007446,
  -4.56523559935519,      -4.65173089980824,      -4.72880744580247,
  -4.79743749076751,      -4.85724052324361,      -4.90844409229379,
  -4.95248457484744,      -4.98903558999084,      -5.01935520927978,
  -5.04389738256082,      -5.06297677321618,      -5.07716591056115,
  -5.08795238885129,      -5.09457802903178,      -5.09646910758147,
  -5.09805117921190,      -5.09323910375321,      -5.08579435904538,
  -5.07580109385102,      -5.05755975890529,      -5.03564993880999,
  -5.00736756957976,      -4.96509673896373,      -4.92310186816408,
  -4.85433590949137,      -4.79291363814269,      -4.68938936781996,
  -4.60668253387820,      -4.45541059237260,      -4.35458956370843,
  -4.14501798325469,      -4.02324984118047,      -3.76696507253240,
  -3.59706560787042,      -3.32857545162272,      -3.07907401636563,
  -2.80915582354951,      -2.50419639837575,      -2.20033587660031,
  -1.88623756749792,      -1.54187737800639,      -1.21814613111141,
 -0.871751094336162,     -0.530254897135803,     -0.197146555849557,
  0.136577164861431,      0.454380148595603,      0.761000151434205,
   1.05131632017050,       1.31949124819132,       1.56741523652175,
   1.79049739805892,       1.98266154375237,       2.14693292913774,
   2.28597342693996,       2.39264122714569,       2.46641825223395,
   2.51471228290353,       2.52649001487208,       2.49464688080853,
   2.44851388159774,       2.39838528163749,       2.33436655077135,
   2.25409992820170,       2.16239258381689,       2.06749613116794,
   1.97479842176582,       1.88561819218097,       1.80820949896022,
   1.74956783886706,       1.70418418830742,       1.67585398062415,
   1.67209464557009,       1.69313184824545,       1.74121786031405,
   1.81717711204739,       1.92129010322954,       2.05387607823807,
   2.21428573935285,       2.40158511037386,       2.61453644547919,
   2.85168017002724,       3.11077744678591,       3.38904948152926,
   3.68413678455739,       3.99247142466248,       4.31183516560780,
   4.63957961513921,       4.97008446943722,       5.30695995168781,
   5.63500167218660,       5.96881162989928,       6.28672856866659,
   6.60090900671800,       6.90472880807607,       7.19281088136067,
   7.47087380401552,       7.73535246020956,       7.98359208903764,
   8.21583740079407,       8.43060479121700,       8.62983142185770,
   8.81643640920844,       8.99051070346617,       9.14968076050637,
   9.29705982134008,       9.43811408186195,       9.56662459418084,
   9.67430571918491,       9.76940693923902,       9.84734960960996,
   9.89554191929840,       9.93936486968965,       9.99280439787169,
   10.0078048229134,       9.96226806398415,       9.91317961573520,
   9.86400214473813,       9.72188511227975,       9.54043438755714,
   9.38489944603994,       9.16534783296569,       9.01727025458012,
   8.78949159959426,       8.28584579406997,       7.93854390914915,
   7.55528012692992,       7.24131651796425,       7.01761461443481,
   6.53953484340049,       6.08603740254494,       5.70706747581750,
   5.26441109863206,       4.82825778041293,       4.45369876702865,
   4.11338633298735,       3.75303173229313,       3.40435451223629,
   3.08698315029473,       2.80260175072035,       2.54708944026464,
   2.31698145579983,       2.11896958316773,       1.94327920206931,
   1.79233856804598,       1.65996154017870,       1.55285192388409,
   1.46777378988845,       1.39037901040042,       1.32883532416728,
   1.27697877262206,       1.21432674176865,       1.14830570011551,
   1.08723958650871,       1.02214218659482,      0.944987850803501,
  0.850530598481662,      0.742448157955449,      0.625221908802865,
  0.489751836406038,      0.329439904055985,      0.150467667980460,
  -2.69098443299436E-002,-0.211973338904167,     -0.385990416613124,
 -0.552771043247399,     -0.705370395871020,     -0.830964447306204,
 -0.918130120743545,      -1.08306350526047,     -0.813442247167167,
  -1.20866845713855,     -0.665340404574263,     -0.799337075481463,
 -0.502003047478292,     -0.628340186640420,      -9.53632873989218E-002,
 -0.128597627409045,      0.292631452445829,      0.235969413573065,
  0.779893537332391,      0.735940049635329,       1.27404762530767,
   1.37669418475712,       1.83814978192687,       2.14406910000102,
   2.60547856270313,       2.96410782308950,       3.39457728602980,
   3.82099418192316,       4.24643132167681,       4.67260459740398,
   5.10767590622106,       5.55410369889172,       5.97292800150418,
   6.34059736008438,       6.71048138901211,       7.08061837004101,
   7.43913349683405,       7.76128797105415,       8.03883367678545,
   8.29931219330208,       8.54771297729456,       8.79809909464291,
   8.96116339412873,       9.10983376424081,       9.35363096770818,
   9.14129033253773,       9.09479954332095,       9.21635856898614,
   9.20691003029131,       9.16091645065158,       9.23972276954451,
   9.18943767529535,       8.89990387232571,       8.77176978190944,
   8.81930863780215,       8.73838651125132,       8.63393494025347,
   8.61203395790562,       8.55122968331386,       8.49079408578536,
   8.43632515671085,       8.42741671396989,       8.44589069482551,
   8.47073937078206,       8.49915484657188,       8.54311503060603,
   8.61290797261590,       8.68452135170458,       8.75053861110366,
   8.83805486146529,       8.94728875493833,       9.02516038371303,
   9.06484019904682,       9.08626325057634,       9.08432534505897,
   9.06254370255456,       8.98251798634018,       8.81980769295451,
   8.64967472346901,       8.49072415460066,       7.63939105349689,
   6.89989571992317,       6.67151123584069,       6.23297746494570,
   4.70564374602921,       4.48461444758391,       3.83341558619055,
   3.00399072387763,       2.12710356314302,       1.50165043714876,
  0.621207434136789,     -0.772862975120267,     -0.957348381249871,
  -2.20198001298990,      -3.05011436818190,      -3.86573074421126,
  -4.78929727445116,      -5.80469037842158,      -6.68185656228296,
  -7.45137413071882,      -8.42505470209597,      -9.13793305776990,
  -10.0052662925040,      -10.7051326094095,      -11.4594069308297,
  -12.1068570644267,      -12.7081047948611,      -13.2774143457626,
  -13.7138049254291,      -14.1644754583250,      -14.4634919444224,
  -14.7593220999530,      -14.9133857058574,      -15.0382187277106,
  -15.0419315126235,      -14.9901738026164,      -14.8371805354244,
  -14.6158082686118,      -14.3058468781334,      -13.9219398413336,
  -13.4606090977760,      -12.9259276797312,      -12.3232454839724,
  -11.6529877011910,      -10.9228534440387,      -10.1330697081775,
  -9.29324532822121,      -8.40354440121031,      -7.47048045563699,
  -6.50241820956604,      -5.50346501219512,      -4.48274285649647,
  -3.43624624385948,      -2.38905820392136,      -1.33642367047722,
 -0.289173967908382,      0.748315900977400,       1.73382252778486,
   2.70007355901374,       3.63030691967745,       4.48186673962542,
   5.25584752002704,       5.96156950202915,       6.56955100078118,
   7.06434435977709,       7.43304916112251,       7.67251243956976,
   7.79966326879873,       7.81054371735532,       7.68808310183721,
   7.44503323201604,       7.10146929608002,       6.66332284670440,
   6.14214573121022,       5.55220341347897,       4.90626546460419,
   4.22469086380833,       3.52544642368524,       2.82145403444239,
   2.12895021926726,       1.46398007873676,      0.840331550812478,
  0.268934132948362,     -0.237978907921587,     -0.675466135317041,
  -1.03282425247745,      -1.31337859187302,      -1.50771031740328,
  -1.62638632787845,      -1.66351479596469,      -1.63252071662317,
  -1.53425880464895,      -1.38148440648380,      -1.18121142611369,
 -0.945210970012627,     -0.683250544086732,     -0.405808657786395,
 -0.122186264522613,      0.159038760526336,      0.430587949755898,
  0.686269459079721,      0.921365153900635,       1.13227407845799,
   1.31694905910953,       1.47459000169248,       1.60555974767556,
   1.71115514754461,       1.79372358531258,       1.85648046166710,
   1.90318954272110,       1.93792892599315,       1.96490882960897,
   1.98841539944117,       2.01266730897658,       2.04147048202241,
   2.07807684661859,       2.12506734963185,       2.18434205897986,
   2.25712972318243,       2.34387315378779,       2.44414392439261,
   2.55677632068255,       2.68008405449131,       2.81195907208257,
   2.94988606054440,       3.09098034874278,       3.23227623866488,
   3.37138782364714,       3.50685057592056,       3.63716904148289,
   3.76025415138737,       3.87518377391334,       3.98293509564728,
   4.08454418294295,       4.17998354790226,       4.26917528841606,
   4.35333999788819,       4.43458811443952,       4.51397022573311,
   4.59141467650580,       4.66835170111963,       4.74630006085218,
   4.82475925489379,       4.90340663435068,       4.98284591145851,
   5.06068400860333,       5.13337787404577,       5.20361251138284,
   5.27158212166067,       5.32473725364969,       5.36330838764898,
   5.39974134044993,       5.42085863099313,       5.41567527847266,
   5.38854419404446,       5.32427668107250,       5.23475419363509,
   5.16348461307841,       5.07650754325165,       4.91446922917897,
   4.73869405051350,       4.59588989638442,       4.43504152484775,
   4.20463289556675,       3.97523110867976,       3.76535688339468,
   3.54438695538454,       3.29142787152686,       3.04764252951938 ;

 time = 1000.0 ;
}
